** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/2x_drive/2bit_comp_2x.sch
**.subckt 2bit_comp_2x L VDD G B1 B0 E A1 A0 VSS
*.iopin VDD
*.ipin B1
*.ipin B0
*.ipin A1
*.iopin VSS
*.ipin A0
*.opin L
*.opin G
*.opin E
x1 VDD B1 net1 A1 VSS my_nxor
x2 VDD B0 net2 A0 VSS my_xor
x3 VDD B0 net2 net3 VSS my_nand
x4 VDD net1 net3 net5 VSS my_nand
x6 VDD B1 net1 net4 VSS my_nor
*  x5 -  my_xor_2x  IS MISSING !!!!
*  x7 -  my_nor_2x  IS MISSING !!!!
*  x8 -  my_nor_2x  IS MISSING !!!!
**.ends

* expanding   symbol:  my_nxor.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nxor.sym
** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nxor.sch
.subckt my_nxor VDD A Out B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin Out
*  M2 -  pfet_03v3  IS MISSING !!!!
*  M4 -  nfet_03v3  IS MISSING !!!!
*  M1 -  pfet_03v3  IS MISSING !!!!
*  M3 -  pfet_03v3  IS MISSING !!!!
*  M5 -  pfet_03v3  IS MISSING !!!!
*  M6 -  nfet_03v3  IS MISSING !!!!
*  M7 -  nfet_03v3  IS MISSING !!!!
*  M8 -  nfet_03v3  IS MISSING !!!!
*  M9 -  pfet_03v3  IS MISSING !!!!
*  M10 -  pfet_03v3  IS MISSING !!!!
*  M11 -  nfet_03v3  IS MISSING !!!!
*  M12 -  nfet_03v3  IS MISSING !!!!
.ends


* expanding   symbol:  my_xor.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_xor.sym
** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_xor.sch
.subckt my_xor VDD A Out B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin Out
*  M2 -  pfet_03v3  IS MISSING !!!!
*  M4 -  nfet_03v3  IS MISSING !!!!
*  M1 -  pfet_03v3  IS MISSING !!!!
*  M3 -  pfet_03v3  IS MISSING !!!!
*  M5 -  pfet_03v3  IS MISSING !!!!
*  M6 -  nfet_03v3  IS MISSING !!!!
*  M7 -  nfet_03v3  IS MISSING !!!!
*  M8 -  nfet_03v3  IS MISSING !!!!
*  M9 -  pfet_03v3  IS MISSING !!!!
*  M10 -  pfet_03v3  IS MISSING !!!!
*  M11 -  nfet_03v3  IS MISSING !!!!
*  M12 -  nfet_03v3  IS MISSING !!!!
.ends


* expanding   symbol:  my_nand.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nand.sym
** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nand.sch
.subckt my_nand VDD A B Out VSS
*.ipin A
*.opin Out
*.ipin B
*.iopin VDD
*.iopin VSS
*  M1 -  nfet_03v3  IS MISSING !!!!
*  M2 -  pfet_03v3  IS MISSING !!!!
*  M3 -  pfet_03v3  IS MISSING !!!!
*  M4 -  nfet_03v3  IS MISSING !!!!
.ends


* expanding   symbol:  my_nor.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nor.sym
** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp4/1x_drive/my_nor.sch
.subckt my_nor VDD A B Out VSS
*.ipin A
*.ipin B
*.iopin VDD
*.iopin VSS
*.opin Out
*  M2 -  pfet_03v3  IS MISSING !!!!
*  M1 -  pfet_03v3  IS MISSING !!!!
*  M3 -  nfet_03v3  IS MISSING !!!!
*  M4 -  nfet_03v3  IS MISSING !!!!
.ends

.end
