magic
tech gf180mcuC
timestamp 1755590146
<< nwell >>
rect 0 63 62 127
<< nmos >>
rect 5 21 11 38
rect 22 21 28 38
rect 33 21 39 38
rect 50 21 56 38
<< pmos >>
rect 19 72 25 106
rect 36 72 42 106
<< ndiff >>
rect -6 32 5 38
rect -6 26 -4 32
rect 2 26 5 32
rect -6 21 5 26
rect 11 29 22 38
rect 11 23 14 29
rect 19 23 22 29
rect 11 21 22 23
rect 28 21 33 38
rect 39 36 50 38
rect 39 23 42 36
rect 47 23 50 36
rect 39 21 50 23
rect 56 32 67 38
rect 56 26 59 32
rect 65 26 67 32
rect 56 21 67 26
<< pdiff >>
rect 9 104 19 106
rect 9 74 11 104
rect 16 74 19 104
rect 9 72 19 74
rect 25 104 36 106
rect 25 79 28 104
rect 33 79 36 104
rect 25 72 36 79
rect 42 104 52 106
rect 42 74 45 104
rect 50 74 52 104
rect 42 72 52 74
<< ndiffc >>
rect -4 26 2 32
rect 14 23 19 29
rect 42 23 47 36
rect 59 26 65 32
<< pdiffc >>
rect 11 74 16 104
rect 28 79 33 104
rect 45 74 50 104
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
<< polysilicon >>
rect 19 106 25 111
rect 36 106 42 111
rect 19 54 25 72
rect 10 52 25 54
rect 10 46 14 52
rect 20 46 25 52
rect 10 44 25 46
rect 5 40 14 44
rect 19 43 25 44
rect 36 67 42 72
rect 36 65 50 67
rect 36 59 42 65
rect 48 59 50 65
rect 36 57 50 59
rect 36 45 42 57
rect 36 43 56 45
rect 19 40 28 43
rect 5 38 11 40
rect 22 38 28 40
rect 33 40 56 43
rect 33 38 39 40
rect 50 38 56 40
rect 5 16 11 21
rect 22 16 28 21
rect 33 16 39 21
rect 50 16 56 21
<< polycontact >>
rect 14 46 20 52
rect 42 59 48 65
<< metal1 >>
rect -6 120 67 127
rect -6 115 11 120
rect 16 115 35 120
rect 40 115 67 120
rect -6 113 67 115
rect 11 104 16 113
rect 28 104 33 106
rect 28 78 33 79
rect 45 104 50 113
rect 11 72 16 74
rect 26 72 28 78
rect 34 72 36 78
rect 45 72 50 74
rect 12 46 14 52
rect 20 46 22 52
rect 28 37 33 72
rect 40 59 42 65
rect 48 59 50 65
rect -5 32 3 34
rect -5 26 -4 32
rect 2 26 3 32
rect -5 24 3 26
rect 14 32 33 37
rect 42 36 47 38
rect 14 29 19 32
rect 14 21 19 23
rect 58 32 66 34
rect 58 26 59 32
rect 65 26 66 32
rect 58 24 66 26
rect 42 14 47 23
rect -6 12 67 14
rect -6 7 11 12
rect 16 7 35 12
rect 40 7 67 12
rect -6 0 67 7
<< via1 >>
rect 28 72 34 78
rect 14 46 20 52
rect 42 59 48 65
rect -4 26 2 32
rect 59 26 65 32
<< metal2 >>
rect 26 78 36 79
rect 26 72 28 78
rect 34 72 36 78
rect 26 71 36 72
rect 40 65 50 66
rect 40 59 42 65
rect 48 59 50 65
rect 40 58 50 59
rect 12 52 22 53
rect 12 46 14 52
rect 20 46 22 52
rect 12 45 22 46
rect -6 32 4 33
rect 57 32 67 33
rect -6 26 -4 32
rect 2 26 59 32
rect 65 26 67 32
rect -6 25 4 26
rect 57 25 67 26
<< labels >>
rlabel metal2 17 49 17 49 1 A
port 1 n
rlabel metal2 45 62 45 62 1 B
port 2 n
rlabel metal2 31 75 31 75 1 Y
port 3 n
rlabel nsubdiffcont 13 118 13 118 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
<< end >>
