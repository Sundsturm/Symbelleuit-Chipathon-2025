magic
tech gf180mcuC
timestamp 1755577130
<< nwell >>
rect -19 63 78 127
<< nmos >>
rect 22 21 28 38
rect 33 21 39 38
<< pmos >>
rect 2 72 8 106
rect 19 72 25 106
rect 36 72 42 106
rect 53 72 59 106
<< ndiff >>
rect 12 29 22 38
rect 12 23 14 29
rect 19 23 22 29
rect 12 21 22 23
rect 28 21 33 38
rect 39 36 49 38
rect 39 23 42 36
rect 47 23 49 36
rect 39 21 49 23
<< pdiff >>
rect -8 104 2 106
rect -8 74 -6 104
rect -1 74 2 104
rect -8 72 2 74
rect 8 104 19 106
rect 8 74 11 104
rect 16 74 19 104
rect 8 72 19 74
rect 25 104 36 106
rect 25 79 28 104
rect 33 79 36 104
rect 25 72 36 79
rect 42 104 53 106
rect 42 74 45 104
rect 50 74 53 104
rect 42 72 53 74
rect 59 104 69 106
rect 59 74 62 104
rect 67 74 69 104
rect 59 72 69 74
<< ndiffc >>
rect 14 23 19 29
rect 42 23 47 36
<< pdiffc >>
rect -6 74 -1 104
rect 11 74 16 104
rect 28 79 33 104
rect 45 74 50 104
rect 62 74 67 104
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
<< polysilicon >>
rect 2 106 8 111
rect 19 106 25 111
rect 36 106 42 111
rect 53 106 59 111
rect 2 54 8 72
rect 19 54 25 72
rect 2 52 25 54
rect 2 48 14 52
rect 11 46 14 48
rect 20 46 25 52
rect 11 44 25 46
rect 19 43 25 44
rect 36 67 42 72
rect 53 67 59 72
rect 36 65 59 67
rect 36 59 42 65
rect 48 61 59 65
rect 48 59 50 61
rect 36 57 50 59
rect 36 43 42 57
rect 19 40 28 43
rect 22 38 28 40
rect 33 40 42 43
rect 33 38 39 40
rect 22 16 28 21
rect 33 16 39 21
<< polycontact >>
rect 14 46 20 52
rect 42 59 48 65
<< metal1 >>
rect -19 120 78 127
rect -19 115 11 120
rect 16 115 35 120
rect 40 115 78 120
rect -19 113 78 115
rect -6 104 -1 106
rect -6 66 -1 74
rect 11 104 16 113
rect 28 104 33 106
rect 28 78 33 79
rect 45 104 50 113
rect 11 72 16 74
rect 26 72 28 78
rect 34 72 36 78
rect 45 72 50 74
rect 62 104 67 106
rect 28 66 33 72
rect -6 61 33 66
rect 28 53 33 61
rect 40 59 42 65
rect 48 59 50 65
rect 62 53 67 74
rect 12 46 14 52
rect 20 46 22 52
rect 28 48 67 53
rect 28 37 33 48
rect 14 32 33 37
rect 42 36 47 38
rect 14 29 19 32
rect 14 21 19 23
rect 42 14 47 23
rect -19 12 78 14
rect -19 7 11 12
rect 16 7 35 12
rect 40 7 78 12
rect -19 0 78 7
<< via1 >>
rect 28 72 34 78
rect 42 59 48 65
rect 14 46 20 52
<< metal2 >>
rect 26 78 36 79
rect 26 72 28 78
rect 34 72 36 78
rect 26 71 36 72
rect 40 65 50 66
rect 40 59 42 65
rect 48 59 50 65
rect 40 58 50 59
rect 12 52 22 53
rect 12 46 14 52
rect 20 46 22 52
rect 12 45 22 46
<< labels >>
rlabel metal2 17 49 17 49 1 A
port 1 n
rlabel metal2 45 62 45 62 1 B
port 2 n
rlabel metal2 31 75 31 75 1 Y
port 3 n
rlabel nsubdiffcont 13 118 13 118 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
<< end >>
