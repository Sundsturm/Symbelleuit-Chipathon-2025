magic
tech gf180mcuD
magscale 1 10
timestamp 1759488065
<< nwell >>
rect -12898 13441 -9740 14153
<< nmos >>
rect -12633 13139 -12573 13309
rect -12465 13139 -12405 13309
rect -12129 13139 -12069 13309
rect -12021 13139 -11961 13309
rect -11685 13139 -11625 13309
rect -11517 13139 -11457 13309
rect -11181 13139 -11121 13309
rect -11013 13139 -10953 13309
rect -10677 13139 -10617 13309
rect -10569 13139 -10509 13309
rect -10233 13139 -10173 13309
rect -10065 13139 -10005 13309
<< pmos >>
rect -12609 13531 -12549 13871
rect -12441 13531 -12381 13871
rect -12105 13531 -12045 13871
rect -11937 13531 -11877 13871
rect -11769 13531 -11709 13871
rect -11601 13531 -11541 13871
rect -11265 13531 -11205 13871
rect -11097 13531 -11037 13871
rect -10761 13531 -10701 13871
rect -10593 13531 -10533 13871
rect -10257 13531 -10197 13871
rect -10089 13531 -10029 13871
<< ndiff >>
rect -12741 13247 -12633 13309
rect -12741 13201 -12710 13247
rect -12664 13201 -12633 13247
rect -12741 13139 -12633 13201
rect -12573 13247 -12465 13309
rect -12573 13201 -12542 13247
rect -12496 13201 -12465 13247
rect -12573 13139 -12465 13201
rect -12405 13247 -12297 13309
rect -12405 13201 -12374 13247
rect -12328 13201 -12297 13247
rect -12405 13139 -12297 13201
rect -12237 13247 -12129 13309
rect -12237 13201 -12206 13247
rect -12160 13201 -12129 13247
rect -12237 13139 -12129 13201
rect -12069 13139 -12021 13309
rect -11961 13247 -11853 13309
rect -11961 13201 -11930 13247
rect -11884 13201 -11853 13247
rect -11961 13139 -11853 13201
rect -11793 13247 -11685 13309
rect -11793 13201 -11762 13247
rect -11716 13201 -11685 13247
rect -11793 13139 -11685 13201
rect -11625 13247 -11517 13309
rect -11625 13201 -11594 13247
rect -11548 13201 -11517 13247
rect -11625 13139 -11517 13201
rect -11457 13247 -11349 13309
rect -11457 13201 -11426 13247
rect -11380 13201 -11349 13247
rect -11457 13139 -11349 13201
rect -11289 13247 -11181 13309
rect -11289 13201 -11258 13247
rect -11212 13201 -11181 13247
rect -11289 13139 -11181 13201
rect -11121 13247 -11013 13309
rect -11121 13201 -11090 13247
rect -11044 13201 -11013 13247
rect -11121 13139 -11013 13201
rect -10953 13247 -10845 13309
rect -10953 13201 -10922 13247
rect -10876 13201 -10845 13247
rect -10953 13139 -10845 13201
rect -10785 13247 -10677 13309
rect -10785 13201 -10754 13247
rect -10708 13201 -10677 13247
rect -10785 13139 -10677 13201
rect -10617 13139 -10569 13309
rect -10509 13247 -10401 13309
rect -10509 13201 -10478 13247
rect -10432 13201 -10401 13247
rect -10509 13139 -10401 13201
rect -10341 13247 -10233 13309
rect -10341 13201 -10310 13247
rect -10264 13201 -10233 13247
rect -10341 13139 -10233 13201
rect -10173 13247 -10065 13309
rect -10173 13201 -10142 13247
rect -10096 13201 -10065 13247
rect -10173 13139 -10065 13201
rect -10005 13247 -9897 13309
rect -10005 13201 -9974 13247
rect -9928 13201 -9897 13247
rect -10005 13139 -9897 13201
<< pdiff >>
rect -12717 13818 -12609 13871
rect -12717 13584 -12686 13818
rect -12640 13584 -12609 13818
rect -12717 13531 -12609 13584
rect -12549 13818 -12441 13871
rect -12549 13584 -12518 13818
rect -12472 13584 -12441 13818
rect -12549 13531 -12441 13584
rect -12381 13818 -12273 13871
rect -12381 13584 -12350 13818
rect -12304 13584 -12273 13818
rect -12381 13531 -12273 13584
rect -12213 13818 -12105 13871
rect -12213 13584 -12182 13818
rect -12136 13584 -12105 13818
rect -12213 13531 -12105 13584
rect -12045 13818 -11937 13871
rect -12045 13584 -12014 13818
rect -11968 13584 -11937 13818
rect -12045 13531 -11937 13584
rect -11877 13818 -11769 13871
rect -11877 13584 -11846 13818
rect -11800 13584 -11769 13818
rect -11877 13531 -11769 13584
rect -11709 13818 -11601 13871
rect -11709 13584 -11678 13818
rect -11632 13584 -11601 13818
rect -11709 13531 -11601 13584
rect -11541 13818 -11433 13871
rect -11541 13584 -11510 13818
rect -11464 13584 -11433 13818
rect -11541 13531 -11433 13584
rect -11373 13818 -11265 13871
rect -11373 13584 -11342 13818
rect -11296 13584 -11265 13818
rect -11373 13531 -11265 13584
rect -11205 13818 -11097 13871
rect -11205 13584 -11174 13818
rect -11128 13584 -11097 13818
rect -11205 13531 -11097 13584
rect -11037 13818 -10929 13871
rect -11037 13584 -11006 13818
rect -10960 13584 -10929 13818
rect -11037 13531 -10929 13584
rect -10869 13818 -10761 13871
rect -10869 13584 -10838 13818
rect -10792 13584 -10761 13818
rect -10869 13531 -10761 13584
rect -10701 13818 -10593 13871
rect -10701 13584 -10670 13818
rect -10624 13584 -10593 13818
rect -10701 13531 -10593 13584
rect -10533 13818 -10425 13871
rect -10533 13584 -10502 13818
rect -10456 13584 -10425 13818
rect -10533 13531 -10425 13584
rect -10365 13818 -10257 13871
rect -10365 13584 -10334 13818
rect -10288 13584 -10257 13818
rect -10365 13531 -10257 13584
rect -10197 13818 -10089 13871
rect -10197 13584 -10166 13818
rect -10120 13584 -10089 13818
rect -10197 13531 -10089 13584
rect -10029 13818 -9921 13871
rect -10029 13584 -9998 13818
rect -9952 13584 -9921 13818
rect -10029 13531 -9921 13584
<< ndiffc >>
rect -12710 13201 -12664 13247
rect -12542 13201 -12496 13247
rect -12374 13201 -12328 13247
rect -12206 13201 -12160 13247
rect -11930 13201 -11884 13247
rect -11762 13201 -11716 13247
rect -11594 13201 -11548 13247
rect -11426 13201 -11380 13247
rect -11258 13201 -11212 13247
rect -11090 13201 -11044 13247
rect -10922 13201 -10876 13247
rect -10754 13201 -10708 13247
rect -10478 13201 -10432 13247
rect -10310 13201 -10264 13247
rect -10142 13201 -10096 13247
rect -9974 13201 -9928 13247
<< pdiffc >>
rect -12686 13584 -12640 13818
rect -12518 13584 -12472 13818
rect -12350 13584 -12304 13818
rect -12182 13584 -12136 13818
rect -12014 13584 -11968 13818
rect -11846 13584 -11800 13818
rect -11678 13584 -11632 13818
rect -11510 13584 -11464 13818
rect -11342 13584 -11296 13818
rect -11174 13584 -11128 13818
rect -11006 13584 -10960 13818
rect -10838 13584 -10792 13818
rect -10670 13584 -10624 13818
rect -10502 13584 -10456 13818
rect -10334 13584 -10288 13818
rect -10166 13584 -10120 13818
rect -9998 13584 -9952 13818
<< psubdiff >>
rect -12834 12955 -12684 12977
rect -12834 12909 -12782 12955
rect -12736 12909 -12684 12955
rect -12834 12887 -12684 12909
rect -12594 12955 -12444 12977
rect -12594 12909 -12542 12955
rect -12496 12909 -12444 12955
rect -12594 12887 -12444 12909
rect -12354 12955 -12204 12977
rect -12354 12909 -12302 12955
rect -12256 12909 -12204 12955
rect -12354 12887 -12204 12909
rect -12114 12955 -11964 12977
rect -12114 12909 -12062 12955
rect -12016 12909 -11964 12955
rect -12114 12887 -11964 12909
rect -11874 12955 -11724 12977
rect -11874 12909 -11822 12955
rect -11776 12909 -11724 12955
rect -11874 12887 -11724 12909
rect -11634 12955 -11484 12977
rect -11634 12909 -11582 12955
rect -11536 12909 -11484 12955
rect -11634 12887 -11484 12909
rect -11394 12955 -11244 12977
rect -11394 12909 -11342 12955
rect -11296 12909 -11244 12955
rect -11394 12887 -11244 12909
rect -11154 12955 -11004 12977
rect -11154 12909 -11102 12955
rect -11056 12909 -11004 12955
rect -11154 12887 -11004 12909
rect -10914 12955 -10764 12977
rect -10914 12909 -10862 12955
rect -10816 12909 -10764 12955
rect -10914 12887 -10764 12909
rect -10674 12955 -10524 12977
rect -10674 12909 -10622 12955
rect -10576 12909 -10524 12955
rect -10674 12887 -10524 12909
rect -10434 12955 -10284 12977
rect -10434 12909 -10382 12955
rect -10336 12909 -10284 12955
rect -10434 12887 -10284 12909
rect -10194 12955 -10044 12977
rect -10194 12909 -10142 12955
rect -10096 12909 -10044 12955
rect -10194 12887 -10044 12909
rect -9954 12955 -9804 12977
rect -9954 12909 -9902 12955
rect -9856 12909 -9804 12955
rect -9954 12887 -9804 12909
<< nsubdiff >>
rect -12834 14099 -12684 14121
rect -12834 14053 -12782 14099
rect -12736 14053 -12684 14099
rect -12834 14031 -12684 14053
rect -12594 14099 -12444 14121
rect -12594 14053 -12542 14099
rect -12496 14053 -12444 14099
rect -12594 14031 -12444 14053
rect -12354 14099 -12204 14121
rect -12354 14053 -12302 14099
rect -12256 14053 -12204 14099
rect -12354 14031 -12204 14053
rect -12114 14099 -11964 14121
rect -12114 14053 -12062 14099
rect -12016 14053 -11964 14099
rect -12114 14031 -11964 14053
rect -11874 14099 -11724 14121
rect -11874 14053 -11822 14099
rect -11776 14053 -11724 14099
rect -11874 14031 -11724 14053
rect -11634 14099 -11484 14121
rect -11634 14053 -11582 14099
rect -11536 14053 -11484 14099
rect -11634 14031 -11484 14053
rect -11394 14099 -11244 14121
rect -11394 14053 -11342 14099
rect -11296 14053 -11244 14099
rect -11394 14031 -11244 14053
rect -11154 14099 -11004 14121
rect -11154 14053 -11102 14099
rect -11056 14053 -11004 14099
rect -11154 14031 -11004 14053
rect -10914 14099 -10764 14121
rect -10914 14053 -10862 14099
rect -10816 14053 -10764 14099
rect -10914 14031 -10764 14053
rect -10674 14099 -10524 14121
rect -10674 14053 -10622 14099
rect -10576 14053 -10524 14099
rect -10674 14031 -10524 14053
rect -10434 14099 -10284 14121
rect -10434 14053 -10382 14099
rect -10336 14053 -10284 14099
rect -10434 14031 -10284 14053
rect -10194 14099 -10044 14121
rect -10194 14053 -10142 14099
rect -10096 14053 -10044 14099
rect -10194 14031 -10044 14053
rect -9954 14099 -9804 14121
rect -9954 14053 -9902 14099
rect -9856 14053 -9804 14099
rect -9954 14031 -9804 14053
<< psubdiffcont >>
rect -12782 12909 -12736 12955
rect -12542 12909 -12496 12955
rect -12302 12909 -12256 12955
rect -12062 12909 -12016 12955
rect -11822 12909 -11776 12955
rect -11582 12909 -11536 12955
rect -11342 12909 -11296 12955
rect -11102 12909 -11056 12955
rect -10862 12909 -10816 12955
rect -10622 12909 -10576 12955
rect -10382 12909 -10336 12955
rect -10142 12909 -10096 12955
rect -9902 12909 -9856 12955
<< nsubdiffcont >>
rect -12782 14053 -12736 14099
rect -12542 14053 -12496 14099
rect -12302 14053 -12256 14099
rect -12062 14053 -12016 14099
rect -11822 14053 -11776 14099
rect -11582 14053 -11536 14099
rect -11342 14053 -11296 14099
rect -11102 14053 -11056 14099
rect -10862 14053 -10816 14099
rect -10622 14053 -10576 14099
rect -10382 14053 -10336 14099
rect -10142 14053 -10096 14099
rect -9902 14053 -9856 14099
<< polysilicon >>
rect -12105 13969 -10197 14009
rect -12609 13871 -12549 13921
rect -12441 13871 -12381 13921
rect -12105 13871 -12045 13969
rect -11937 13871 -11877 13921
rect -11769 13871 -11709 13921
rect -11601 13871 -11541 13921
rect -11265 13871 -11205 13969
rect -11097 13871 -11037 13921
rect -10761 13871 -10701 13921
rect -10593 13871 -10533 13921
rect -10257 13871 -10197 13969
rect -10089 13871 -10029 13921
rect -12609 13503 -12549 13531
rect -12633 13455 -12549 13503
rect -12633 13409 -12614 13455
rect -12568 13409 -12549 13455
rect -12633 13379 -12549 13409
rect -12633 13309 -12573 13379
rect -12441 13377 -12381 13531
rect -12105 13511 -12045 13531
rect -12129 13471 -12045 13511
rect -12465 13337 -12381 13377
rect -12169 13447 -12069 13471
rect -12169 13401 -12150 13447
rect -12104 13401 -12069 13447
rect -12169 13371 -12069 13401
rect -11937 13462 -11877 13531
rect -11769 13462 -11709 13531
rect -11601 13503 -11541 13531
rect -11601 13463 -11457 13503
rect -11937 13441 -11709 13462
rect -11937 13395 -11843 13441
rect -11797 13395 -11709 13441
rect -11937 13377 -11709 13395
rect -12465 13309 -12405 13337
rect -12129 13309 -12069 13371
rect -12021 13337 -11625 13377
rect -12021 13309 -11961 13337
rect -11685 13309 -11625 13337
rect -11517 13309 -11457 13463
rect -11265 13377 -11205 13531
rect -11097 13503 -11037 13531
rect -10761 13503 -10701 13531
rect -11097 13463 -10701 13503
rect -10593 13511 -10533 13531
rect -10593 13471 -10509 13511
rect -10822 13441 -10723 13463
rect -10822 13395 -10795 13441
rect -10749 13395 -10723 13441
rect -10822 13377 -10723 13395
rect -10569 13447 -10469 13471
rect -10569 13401 -10550 13447
rect -10504 13401 -10469 13447
rect -11265 13337 -11121 13377
rect -11181 13309 -11121 13337
rect -11013 13337 -10617 13377
rect -11013 13309 -10953 13337
rect -10677 13309 -10617 13337
rect -10569 13371 -10469 13401
rect -10257 13377 -10197 13531
rect -10089 13503 -10029 13531
rect -10089 13455 -10005 13503
rect -10089 13409 -10070 13455
rect -10024 13409 -10005 13455
rect -10089 13379 -10005 13409
rect -10569 13309 -10509 13371
rect -10257 13337 -10173 13377
rect -10233 13309 -10173 13337
rect -10065 13309 -10005 13379
rect -12633 13089 -12573 13139
rect -12465 13041 -12405 13139
rect -12129 13089 -12069 13139
rect -12021 13089 -11961 13139
rect -11685 13089 -11625 13139
rect -11517 13041 -11457 13139
rect -11181 13089 -11121 13139
rect -11013 13089 -10953 13139
rect -10677 13089 -10617 13139
rect -10569 13041 -10509 13139
rect -10233 13089 -10173 13139
rect -10065 13089 -10005 13139
rect -12465 13001 -10509 13041
<< polycontact >>
rect -12614 13409 -12568 13455
rect -12150 13401 -12104 13447
rect -11843 13395 -11797 13441
rect -10795 13395 -10749 13441
rect -10550 13401 -10504 13447
rect -10070 13409 -10024 13455
<< metal1 >>
rect -12898 14099 -9740 14153
rect -12898 14053 -12782 14099
rect -12736 14053 -12542 14099
rect -12496 14053 -12302 14099
rect -12256 14053 -12062 14099
rect -12016 14053 -11822 14099
rect -11776 14053 -11582 14099
rect -11536 14053 -11342 14099
rect -11296 14053 -11102 14099
rect -11056 14053 -10862 14099
rect -10816 14053 -10622 14099
rect -10576 14053 -10382 14099
rect -10336 14053 -10142 14099
rect -10096 14053 -9902 14099
rect -9856 14053 -9740 14099
rect -12898 14013 -9740 14053
rect -12690 13818 -12638 13871
rect -12690 13584 -12686 13818
rect -12640 13584 -12638 13818
rect -12690 13583 -12638 13584
rect -12743 13531 -12638 13583
rect -12521 13818 -12469 14013
rect -12521 13584 -12518 13818
rect -12472 13584 -12469 13818
rect -12521 13531 -12469 13584
rect -12354 13818 -12302 13874
rect -12354 13584 -12350 13818
rect -12304 13584 -12302 13818
rect -12743 13462 -12691 13531
rect -12354 13513 -12302 13584
rect -12185 13818 -12133 14013
rect -12185 13584 -12182 13818
rect -12136 13584 -12133 13818
rect -12185 13559 -12133 13584
rect -12017 13818 -11965 13871
rect -12017 13584 -12014 13818
rect -11968 13584 -11965 13818
rect -12792 13412 -12691 13462
rect -12792 13360 -12768 13412
rect -12716 13360 -12691 13412
rect -12633 13458 -12549 13475
rect -12633 13406 -12617 13458
rect -12565 13406 -12549 13458
rect -12633 13379 -12549 13406
rect -12378 13471 -12302 13513
rect -12378 13419 -12367 13471
rect -12315 13419 -12302 13471
rect -12792 13309 -12691 13360
rect -12378 13337 -12302 13419
rect -12169 13485 -12069 13511
rect -12169 13433 -12153 13485
rect -12101 13433 -12069 13485
rect -12169 13401 -12150 13433
rect -12104 13401 -12069 13433
rect -12169 13371 -12069 13401
rect -12743 13257 -12661 13309
rect -12713 13247 -12661 13257
rect -12713 13201 -12710 13247
rect -12664 13201 -12661 13247
rect -12713 13134 -12661 13201
rect -12545 13247 -12493 13309
rect -12545 13201 -12542 13247
rect -12496 13201 -12493 13247
rect -12545 13023 -12493 13201
rect -12378 13247 -12326 13337
rect -12017 13309 -11965 13584
rect -11849 13818 -11797 14013
rect -11849 13584 -11846 13818
rect -11800 13584 -11797 13818
rect -11849 13531 -11797 13584
rect -11681 13818 -11629 13878
rect -11681 13584 -11678 13818
rect -11632 13584 -11629 13818
rect -11681 13512 -11629 13584
rect -11541 13818 -11433 13871
rect -11541 13779 -11510 13818
rect -11464 13779 -11433 13818
rect -11541 13623 -11513 13779
rect -11461 13623 -11433 13779
rect -11541 13584 -11510 13623
rect -11464 13584 -11433 13623
rect -11541 13560 -11433 13584
rect -11345 13818 -11293 14013
rect -11345 13584 -11342 13818
rect -11296 13584 -11293 13818
rect -11345 13560 -11293 13584
rect -11177 13818 -11125 13871
rect -11177 13584 -11174 13818
rect -11128 13584 -11125 13818
rect -11177 13512 -11125 13584
rect -11037 13818 -10929 13871
rect -11037 13779 -11006 13818
rect -10960 13779 -10929 13818
rect -11037 13623 -11009 13779
rect -10957 13623 -10929 13779
rect -11037 13584 -11006 13623
rect -10960 13584 -10929 13623
rect -11037 13560 -10929 13584
rect -10841 13818 -10789 14013
rect -10841 13584 -10838 13818
rect -10792 13584 -10789 13818
rect -10841 13531 -10789 13584
rect -10673 13818 -10621 13871
rect -10673 13584 -10670 13818
rect -10624 13584 -10621 13818
rect -11902 13444 -11745 13462
rect -11681 13460 -11125 13512
rect -11902 13392 -11846 13444
rect -11794 13392 -11745 13444
rect -10822 13444 -10723 13463
rect -11902 13377 -11745 13392
rect -11429 13357 -10873 13409
rect -10822 13392 -10798 13444
rect -10746 13392 -10723 13444
rect -10822 13377 -10723 13392
rect -12378 13201 -12374 13247
rect -12328 13201 -12326 13247
rect -12378 13139 -12326 13201
rect -12209 13247 -12157 13309
rect -12209 13201 -12206 13247
rect -12160 13201 -12157 13247
rect -12209 13023 -12157 13201
rect -12021 13247 -11853 13309
rect -12021 13219 -11930 13247
rect -11884 13219 -11853 13247
rect -12021 13167 -11933 13219
rect -11881 13167 -11853 13219
rect -12021 13139 -11853 13167
rect -11766 13247 -11714 13309
rect -11766 13201 -11762 13247
rect -11716 13201 -11714 13247
rect -11766 13123 -11714 13201
rect -11625 13251 -11517 13285
rect -11625 13199 -11597 13251
rect -11545 13199 -11517 13251
rect -11625 13171 -11517 13199
rect -11429 13247 -11377 13357
rect -11429 13201 -11426 13247
rect -11380 13201 -11377 13247
rect -11429 13171 -11377 13201
rect -11261 13247 -11209 13309
rect -11261 13201 -11258 13247
rect -11212 13201 -11209 13247
rect -11261 13123 -11209 13201
rect -11766 13071 -11209 13123
rect -11094 13247 -11042 13309
rect -11094 13201 -11090 13247
rect -11044 13201 -11042 13247
rect -11094 13023 -11042 13201
rect -10925 13247 -10873 13357
rect -10673 13309 -10621 13584
rect -10505 13818 -10453 14013
rect -10505 13584 -10502 13818
rect -10456 13584 -10453 13818
rect -10505 13559 -10453 13584
rect -10337 13818 -10285 13874
rect -10337 13584 -10334 13818
rect -10288 13584 -10285 13818
rect -10337 13513 -10285 13584
rect -10169 13818 -10117 14013
rect -10169 13584 -10166 13818
rect -10120 13584 -10117 13818
rect -10169 13531 -10117 13584
rect -10001 13818 -9949 13871
rect -10001 13584 -9998 13818
rect -9952 13584 -9949 13818
rect -10001 13583 -9949 13584
rect -10001 13531 -9897 13583
rect -10569 13485 -10469 13511
rect -10569 13433 -10553 13485
rect -10501 13433 -10469 13485
rect -10569 13401 -10550 13433
rect -10504 13401 -10469 13433
rect -10569 13371 -10469 13401
rect -10337 13471 -10261 13513
rect -10337 13419 -10324 13471
rect -10272 13419 -10261 13471
rect -10337 13377 -10261 13419
rect -10089 13458 -10005 13480
rect -10089 13406 -10073 13458
rect -10021 13406 -10005 13458
rect -10089 13379 -10005 13406
rect -9949 13462 -9897 13531
rect -9949 13412 -9846 13462
rect -10925 13201 -10922 13247
rect -10876 13201 -10873 13247
rect -10925 13139 -10873 13201
rect -10785 13247 -10617 13309
rect -10785 13219 -10754 13247
rect -10708 13219 -10617 13247
rect -10785 13167 -10757 13219
rect -10705 13167 -10617 13219
rect -10785 13139 -10617 13167
rect -10481 13247 -10429 13309
rect -10481 13201 -10478 13247
rect -10432 13201 -10429 13247
rect -10481 13023 -10429 13201
rect -10313 13247 -10261 13377
rect -9949 13360 -9921 13412
rect -9869 13360 -9846 13412
rect -9949 13309 -9846 13360
rect -10313 13201 -10310 13247
rect -10264 13201 -10261 13247
rect -10313 13139 -10261 13201
rect -10145 13247 -10093 13309
rect -10145 13201 -10142 13247
rect -10096 13201 -10093 13247
rect -10145 13023 -10093 13201
rect -9977 13257 -9897 13309
rect -9977 13247 -9925 13257
rect -9977 13201 -9974 13247
rect -9928 13201 -9925 13247
rect -9977 13140 -9925 13201
rect -12862 12955 -9776 13023
rect -12862 12909 -12782 12955
rect -12736 12909 -12542 12955
rect -12496 12909 -12302 12955
rect -12256 12909 -12062 12955
rect -12016 12909 -11822 12955
rect -11776 12909 -11582 12955
rect -11536 12909 -11342 12955
rect -11296 12909 -11102 12955
rect -11056 12909 -10862 12955
rect -10816 12909 -10622 12955
rect -10576 12909 -10382 12955
rect -10336 12909 -10142 12955
rect -10096 12909 -9902 12955
rect -9856 12909 -9776 12955
rect -12862 12883 -9776 12909
<< via1 >>
rect -12768 13360 -12716 13412
rect -12617 13455 -12565 13458
rect -12617 13409 -12614 13455
rect -12614 13409 -12568 13455
rect -12568 13409 -12565 13455
rect -12617 13406 -12565 13409
rect -12367 13419 -12315 13471
rect -12153 13447 -12101 13485
rect -12153 13433 -12150 13447
rect -12150 13433 -12104 13447
rect -12104 13433 -12101 13447
rect -11513 13623 -11510 13779
rect -11510 13623 -11464 13779
rect -11464 13623 -11461 13779
rect -11009 13623 -11006 13779
rect -11006 13623 -10960 13779
rect -10960 13623 -10957 13779
rect -11846 13441 -11794 13444
rect -11846 13395 -11843 13441
rect -11843 13395 -11797 13441
rect -11797 13395 -11794 13441
rect -11846 13392 -11794 13395
rect -10798 13441 -10746 13444
rect -10798 13395 -10795 13441
rect -10795 13395 -10749 13441
rect -10749 13395 -10746 13441
rect -10798 13392 -10746 13395
rect -11933 13201 -11930 13219
rect -11930 13201 -11884 13219
rect -11884 13201 -11881 13219
rect -11933 13167 -11881 13201
rect -11597 13247 -11545 13251
rect -11597 13201 -11594 13247
rect -11594 13201 -11548 13247
rect -11548 13201 -11545 13247
rect -11597 13199 -11545 13201
rect -10553 13447 -10501 13485
rect -10553 13433 -10550 13447
rect -10550 13433 -10504 13447
rect -10504 13433 -10501 13447
rect -10324 13419 -10272 13471
rect -10073 13455 -10021 13458
rect -10073 13409 -10070 13455
rect -10070 13409 -10024 13455
rect -10024 13409 -10021 13455
rect -10073 13406 -10021 13409
rect -10757 13201 -10754 13219
rect -10754 13201 -10708 13219
rect -10708 13201 -10705 13219
rect -10757 13167 -10705 13201
rect -9921 13360 -9869 13412
<< metal2 >>
rect -11601 13779 -11433 13871
rect -11601 13623 -11513 13779
rect -11461 13730 -11433 13779
rect -11037 13779 -10929 13871
rect -11037 13730 -11009 13779
rect -11461 13670 -11009 13730
rect -11461 13623 -11433 13670
rect -11601 13560 -11433 13623
rect -11037 13623 -11009 13670
rect -10957 13623 -10929 13779
rect -11037 13560 -10929 13623
rect -12633 13475 -12573 13503
rect -12792 13412 -12693 13462
rect -12792 13360 -12768 13412
rect -12716 13360 -12693 13412
rect -12792 13309 -12693 13360
rect -12633 13458 -12549 13475
rect -12633 13406 -12617 13458
rect -12565 13406 -12549 13458
rect -12633 13379 -12549 13406
rect -12378 13471 -12302 13513
rect -12378 13419 -12367 13471
rect -12315 13419 -12302 13471
rect -12633 13139 -12573 13379
rect -12378 13357 -12302 13419
rect -12169 13485 -12085 13511
rect -12169 13433 -12153 13485
rect -12101 13433 -12085 13485
rect -12169 13417 -12085 13433
rect -11937 13444 -11709 13462
rect -11937 13392 -11846 13444
rect -11794 13392 -11709 13444
rect -11937 13377 -11709 13392
rect -11937 13357 -11877 13377
rect -12378 13337 -11877 13357
rect -12362 13297 -11877 13337
rect -11601 13285 -11541 13560
rect -10569 13485 -10485 13511
rect -10822 13444 -10723 13463
rect -10822 13392 -10798 13444
rect -10746 13392 -10723 13444
rect -10569 13433 -10553 13485
rect -10501 13433 -10485 13485
rect -10569 13417 -10485 13433
rect -10337 13471 -10261 13513
rect -10065 13480 -10005 13503
rect -10337 13419 -10324 13471
rect -10272 13419 -10261 13471
rect -10822 13377 -10723 13392
rect -10783 13357 -10723 13377
rect -10337 13377 -10261 13419
rect -10089 13458 -10005 13480
rect -10089 13406 -10073 13458
rect -10021 13406 -10005 13458
rect -10089 13379 -10005 13406
rect -10337 13357 -10277 13377
rect -10783 13297 -10277 13357
rect -11625 13251 -11517 13285
rect -12021 13219 -11853 13235
rect -12021 13167 -11933 13219
rect -11881 13167 -11853 13219
rect -11625 13199 -11597 13251
rect -11545 13199 -11517 13251
rect -11625 13171 -11517 13199
rect -10785 13219 -10617 13235
rect -12021 13139 -11853 13167
rect -11601 13152 -11541 13171
rect -10785 13167 -10757 13219
rect -10705 13167 -10617 13219
rect -12633 13079 -11853 13139
rect -10785 13139 -10617 13167
rect -10065 13139 -10005 13379
rect -9945 13412 -9846 13462
rect -9945 13360 -9921 13412
rect -9869 13360 -9846 13412
rect -9945 13309 -9846 13360
rect -10785 13079 -10005 13139
<< labels >>
flabel metal2 s -12128 13463 -12128 13463 2 FreeSans 448 0 0 0 B
port 1 nsew
flabel metal2 s -10530 13464 -10530 13464 2 FreeSans 448 0 0 0 A
port 2 nsew
flabel metal2 s -12768 13343 -12768 13343 2 FreeSans 700 0 0 0 L
port 3 nsew
flabel metal2 s -11586 13378 -11586 13378 2 FreeSans 700 0 0 0 E
port 4 nsew
flabel metal2 s -9881 13336 -9881 13336 2 FreeSans 700 0 0 0 G
port 5 nsew
flabel metal1 s -10244 14085 -10244 14085 2 FreeSans 576 0 0 0 VDD
port 6 nsew
flabel metal1 s -10244 12936 -10244 12936 2 FreeSans 576 0 0 0 VSS
port 7 nsew
<< properties >>
string path -61.660 66.950 -61.660 66.635 -59.535 66.635 -59.535 67.160 
<< end >>
