* NGSPICE file created from gf180mcu_gp9t3v3__comp2_2.ext - technology: gf180mcuD

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

.subckt gf180mcu_gp9t3v3__comp2_2 B A G L E VDD VSS
X0 VDD a_n12969_13089# L VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X1 G a_n10617_13139# VSS VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.2295p ps=1.39u w=0.85u l=0.3u
X2 VSS B a_n11961_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X3 VDD A a_n10617_13139# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X4 L a_n12969_13089# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X5 a_n12573_13139# A VDD VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X6 a_n11877_13531# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X7 a_n12573_13139# A VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X8 VSS a_n11013_13089# a_n11625_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X9 VSS a_n10617_13139# G VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X10 a_n11625_13139# a_n11013_13089# VSS VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.2295p ps=1.39u w=0.85u l=0.3u
X11 a_n10449_13139# a_n11013_13089# a_n10617_13139# VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X12 VDD B a_n11877_13531# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X13 VDD a_n10617_13139# G VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X14 VSS a_n12969_13089# L VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.2295p ps=1.39u w=0.85u l=0.3u
X15 L a_n12969_13089# VSS VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X16 a_n11625_13139# A E VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.2295p ps=1.39u w=0.85u l=0.3u
X17 VSS B a_n11013_13089# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X18 E a_n11013_13089# a_n11877_13531# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X19 G a_n10617_13139# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X20 E a_n12573_13139# a_n11961_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X21 E A a_n11625_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X22 a_n11877_13531# A E VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X23 a_n12969_13089# a_n12573_13139# a_n12237_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X24 a_n12969_13089# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X25 E A a_n11877_13531# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X26 VSS A a_n10449_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X27 a_n11877_13531# a_n12573_13139# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X28 VDD a_n12573_13139# a_n12969_13089# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X29 VDD B a_n11013_13089# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X30 a_n12237_13139# B VSS VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X31 a_n10617_13139# a_n11013_13089# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
.ends

