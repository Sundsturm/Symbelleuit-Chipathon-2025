  X � 	   0 � 	   0  LIB  >A�7KƧ�9D�/��ZT � 	   0 � 	   0  gf180mcu_gp9t3v3__comp2_1         ,��� ���� m��A m��A ���� �          ,��
 )��
 ���� ���� )��
 )          ,��� )��� ���� ���� )��� )          ,��f )��f ���T ���T )��f )          ,�� )�� ��� ��� )�� )          ,��� )��� ���� ���� )��� )          ,��!v )��!v ���$d ���$d )��!v )          ,��&& )��&& ���) ���) )��&& )          ,��*� )��*� ���-� ���-� )��*� )          ,��/� )��/� ���2t ���2t )��/� )          ,��46 )��46 ���7$ ���7$ )��46 )          ,��8� )��8� ���;� ���;� )��8� )          ,��� G��� ���K ���K G��� G          ,��w G��w ��� � ��� � G��w G          ,��!� G��!� ���*� ���*� G��!� G          ,��+� G��+� ���4c ���4c G��+� G          ,��5� G��5� ���>; ���>; G��5� G          ,��'  ���' ���� ����  ���'  �          ,���  ���� ��� ���  ����  �          ,���  ���� ���"W ���"W  ����  �          ,��#�  ���#� ���,/ ���,/  ���#�  �          ,��-[  ���-[ ���4� ���4�  ���-[  �          ,��6  ���6 ���>� ���>�  ���6  �          ,��
  ����
  �a���  �a���  ����
  ��          ,���  �����  �a���  �a���  �����  ��          ,��f  ����f  �a��T  �a��T  ����f  ��          ,��  ����  �a��  �a��  ����  ��          ,���  �����  �a���  �a���  �����  ��          ,��!v  ����!v  �a��$d  �a��$d  ����!v  ��          ,��&&  ����&&  �a��)  �a��)  ����&&  ��          ,��*�  ����*�  �a��-�  �a��-�  ����*�  ��          ,��/�  ����/�  �a��2t  �a��2t  ����/�  ��          ,��46  ����46  �a��7$  �a��7$  ����46  ��          ,��8�  ����8�  �a��;�  �a��;�  ����8�  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��V )��V ���D ���D )��V )          ,��=� )��=� ���@� ���@� )��=� )          ,��
 )��
 ���� ���� )��
 )          ,��
 )��
 ���� ���� )��
 )          ,��=� )��=� ���@� ���@� )��=� )          ,��V )��V ���D ���D )��V )          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��8�  ����8�  �a��;�  �a��;�  ����8�  ��          ,��46  ����46  �a��7$  �a��7$  ����46  ��          ,��/�  ����/�  �a��2t  �a��2t  ����/�  ��          ,��*�  ����*�  �a��-�  �a��-�  ����*�  ��          ,��&&  ����&&  �a��)  �a��)  ����&&  ��          ,��!v  ����!v  �a��$d  �a��$d  ����!v  ��          ,���  �����  �a���  �a���  �����  ��          ,��  ����  �a��  �a��  ����  ��          ,��f  ����f  �a��T  �a��T  ����f  ��          ,���  �����  �a���  �a���  �����  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��6  ���6 ���>� ���>�  ���6  �          ,��-[  ���-[ ���4� ���4�  ���-[  �          ,��#�  ���#� ���,/ ���,/  ���#�  �          ,���  ���� ���"W ���"W  ����  �          ,���  ���� ��� ���  ����  �          ,��'  ���' ���� ����  ���'  �          ,��5� G��5� ���>; ���>; G��5� G          ,��+� G��+� ���4c ���4c G��+� G          ,��!� G��!� ���*� ���*� G��!� G          ,��w G��w ��� � ��� � G��w G          ,��� G��� ���K ���K G��� G          ,��8� )��8� ���;� ���;� )��8� )          ,��46 )��46 ���7$ ���7$ )��46 )          ,��/� )��/� ���2t ���2t )��/� )          ,��*� )��*� ���-� ���-� )��*� )          ,��&& )��&& ���) ���) )��&& )          ,��!v )��!v ���$d ���$d )��!v )          ,��� )��� ���� ���� )��� )          ,�� )�� ��� ��� )�� )          ,��f )��f ���T ���T )��f )          ,��� )��� ���� ���� )��� )          ,��
 )��
 ���� ���� )��
 )           ,��V ��V m��@� m��@� ��V            ,��	� ��	� �� �� ��	�            ,��� ��� ��� ��� ���            ,��R ��R ��h ��h ��R            ,�� �� �� �� ��            ,��� ��� ��� ��� ���            ,��!b ��!b ��$x ��$x ��!b            ,��& ��& ��)( ��)( ��&            ,��*� ��*� ��-� ��-� ��*�            ,��/r ��/r ��2� ��2� ��/r            ,��4" ��4" ��78 ��78 ��4"            ,��8� ��8� ��;� ��;� ��8�            ,��] ���] ���� ���� ���] �           ,��5 ���5 ���I ���I ���5 �           ,��� ���� ���!! ���!! ���� �           ,��$� ���$� ���*� ���*� ���$� �           ,��.� ���.� ���3� ���3� ���.� �           ,��7= ���7= ���=} ���=} ���7= �           ,���  ����� ���?S ���?S  �����  ��           ,��]  ����]  �����  �����  ����]  ��           ,��5  ����5  ����I  ����I  ����5  ��           ,���  �����  ����!!  ����!!  �����  ��           ,��$�  ����$�  ����*�  ����*�  ����$�  ��           ,��.�  ����.�  ����3�  ����3�  ����.�  ��           ,��7=  ����7=  ����=}  ����=}  ����7=  ��           ,��V ��V ��X ��X ��V            ,��=� ��=� ��@� ��@� ��=�            ,��	� ��	� �� �� ��	�            ,��	� ��	� �� �� ��	�            ,��=� ��=� ��@� ��@� ��=�            ,��V ��V ��X ��X ��V            ,��7=  ����7=  ����=}  ����=}  ����7=  ��           ,��.�  ����.�  ����3�  ����3�  ����.�  ��           ,��$�  ����$�  ����*�  ����*�  ����$�  ��           ,���  �����  ����!!  ����!!  �����  ��           ,��5  ����5  ����I  ����I  ����5  ��           ,��]  ����]  �����  �����  ����]  ��           ,���  ����� ���?S ���?S  �����  ��           ,��7= ���7= ���=} ���=} ���7= �           ,��.� ���.� ���3� ���3� ���.� �           ,��$� ���$� ���*� ���*� ���$� �           ,��� ���� ���!! ���!! ���� �           ,��5 ���5 ���I ���I ���5 �           ,��] ���] ���� ���� ���] �           ,��8� ��8� ��;� ��;� ��8�            ,��4" ��4" ��78 ��78 ��4"            ,��/r ��/r ��2� ��2� ��/r            ,��*� ��*� ��-� ��-� ��*�            ,��& ��& ��)( ��)( ��&            ,��!b ��!b ��$x ��$x ��!b            ,��� ��� ��� ��� ���            ,�� �� �� �� ��            ,��R ��R ��h ��h ��R            ,��� ��� ��� ��� ���            ,��	� ��	� �� �� ��	�            ,��V ��V m��@� m��@� ��V           ,��� ���� ��� ��� ���� �          ,��� ���� ���} ���} ���� �          ,��# ���# ���)U ���)U ���# �          ,��,� ���,� ���3- ���3- ���,� �          ,��6� ���6� ���= ���= ���6� �          ,��� ���� ���>� ���>� ���� �          ,��� a��� ��� ��� a��� a          ,��� a��� ���} ���} a��� a          ,��# a��# ���)U ���)U a��# a          ,��,� a��,� ���3- ���3- a��,� a          ,��6� a��6� ���= ���= a��6� a          ,���  �����  �u���  �u���  �����  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��R  ����R  �u��h  �u��h  ����R  ��          ,��  ����  �u��  �u��  ����  ��          ,���  �����  �u���  �u���  �����  ��          ,��!b  ����!b  �u��$x  �u��$x  ����!b  ��          ,��&  ����&  �u��)(  �u��)(  ����&  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��          ,��/r  ����/r  �u��2�  �u��2�  ����/r  ��          ,��4"  ����4"  �u��78  �u��78  ����4"  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��	�  ����	�  �u��  �u��  ����	�  ��          ,��B  ����B  �u��X  �u��X  ����B  ��          ,��B  ����B  �u��X  �u��X  ����B  ��          ,��	�  ����	�  �u��  �u��  ����	�  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��4"  ����4"  �u��78  �u��78  ����4"  ��          ,��/r  ����/r  �u��2�  �u��2�  ����/r  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��          ,��&  ����&  �u��)(  �u��)(  ����&  ��          ,��!b  ����!b  �u��$x  �u��$x  ����!b  ��          ,���  �����  �u���  �u���  �����  ��          ,��  ����  �u��  �u��  ����  ��          ,��R  ����R  �u��h  �u��h  ����R  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,���  �����  �u���  �u���  �����  ��          ,��6� a��6� ���= ���= a��6� a          ,��,� a��,� ���3- ���3- a��,� a          ,��# a��# ���)U ���)U a��# a          ,��� a��� ���} ���} a��� a          ,��� a��� ��� ��� a��� a          ,��� ���� ���>� ���>� ���� �          ,��6� ���6� ���= ���= ���6� �          ,��,� ���,� ���3- ���3- ���,� �          ,��# ���# ���)U ���)U ���# �          ,��� ���� ���} ���} ���� �          ,��� ���� ��� ��� ���� �          ,��� ���� ���8� ���8� ���� �          ,��	� ���	� ���
� ���
� ���	� �          ,��	C O��	C ���
� ���
� O��	C O          ,��	C  ����	C O��
o O��
o  ����	C  ��          ,�� E�� ���/ ���/ E�� E          ,��� ���� ���� ���� ���� �          ,��� }��� E��/ E��/ }��� }          ,�� ��� ���� ���� ��� �          ,���  ����� }��� }���  �����  ��          ,��  ���� ���G ���G  ����  ��          ,��� ���� ��� ��� ���� �          ,��# ���# ���O ���O ���# �          ,��k ���k ���� ���� ���k �          ,��k ���k ��� ; ��� ; ���k �          ,��� E��� ���O ���O E��� E          ,��7 }��7 E��� E��� }��7 }          ,��7  ����7 }��c }��c  ����7  ��          ,���  ����� }��� }���  �����  ��          ,��  ���� ��� ; ��� ;  ����  ��          ,��#� E��#� ���%' ���%' E��#� E          ,��'C ���'C ���(o ���(o ���'C �          ,��-� ���-� ���.� ���.� ���-� �          ,��'C ���'C ���.� ���.� ���'C �          ,��1 ���1 ���2G ���2G ���1 �          ,��1 ���1 ���2� ���2� ���1 �          ,��,� E��,� ���.� ���.� E��,� E          ,��#� }��#� E��&� E��&� }��#� }          ,��%�  ����%� }��&� }��&�  ����%�  ��          ,��(� }��(� E��0� E��0� }��(� }          ,��(�  ����(� }��* }��*  ����(�  ��          ,��/w  ����/w }��0� }��0�  ����/w  ��          ,��1�  ����1� ���2� ���2�  ����1�  ��          ,��7� E��7� ���8� ���8� E��7� E          ,��:� ���:� ���< ���< ���:� �          ,��:� O��:� ���<� ���<� O��:� O          ,��7� }��7� E��9O E��9O }��7� }          ,��8#  ����8# }��9O }��9O  ����8#  ��          ,��;k  ����;k O��<� O��<�  ����;k  ��          ,���  �����  ����2�  ����2�  �����  ��          ,���  �����  ����2�  ����2�  �����  ��          ,��;k  ����;k O��<� O��<�  ����;k  ��          ,��8#  ����8# }��9O }��9O  ����8#  ��          ,��7� }��7� E��9O E��9O }��7� }          ,��:� O��:� ���<� ���<� O��:� O          ,��:� ���:� ���< ���< ���:� �          ,��7� E��7� ���8� ���8� E��7� E          ,��1�  ����1� ���2� ���2�  ����1�  ��          ,��/w  ����/w }��0� }��0�  ����/w  ��          ,��(�  ����(� }��* }��*  ����(�  ��          ,��(� }��(� E��0� E��0� }��(� }          ,��%�  ����%� }��&� }��&�  ����%�  ��          ,��#� }��#� E��&� E��&� }��#� }          ,��,� E��,� ���.� ���.� E��,� E          ,��1 ���1 ���2� ���2� ���1 �          ,��1 ���1 ���2G ���2G ���1 �          ,��'C ���'C ���.� ���.� ���'C �          ,��-� ���-� ���.� ���.� ���-� �          ,��'C ���'C ���(o ���(o ���'C �          ,��#� E��#� ���%' ���%' E��#� E          ,��  ���� ��� ; ��� ;  ����  ��          ,���  ����� }��� }���  �����  ��          ,��7  ����7 }��c }��c  ����7  ��          ,��7 }��7 E��� E��� }��7 }          ,��� E��� ���O ���O E��� E          ,��k ���k ��� ; ��� ; ���k �          ,��k ���k ���� ���� ���k �          ,��# ���# ���O ���O ���# �          ,��� ���� ��� ��� ���� �          ,��  ���� ���G ���G  ����  ��          ,���  ����� }��� }���  �����  ��          ,�� ��� ���� ���� ��� �          ,��� }��� E��/ E��/ }��� }          ,��� ���� ���� ���� ���� �          ,�� E�� ���/ ���/ E�� E          ,��	C  ����	C O��
o O��
o  ����	C  ��          ,��	C O��	C ���
� ���
� O��	C O          ,��	� ���	� ���
� ���
� ���	� �          ,��� ���� ���8� ���8� ���� �      !    ,��" ���" x��#[ x��#[ ���" �      !    ,��" ��" ���#[ ���#[ ��"       !    ,��" +��" ��#[ ��#[ +��" +      !    ,��" 	U��" 
1��#[ 
1��#[ 	U��" 	U      !    ,��"  ���"  ����#[  ����#[  ���"  �      !    ,��"  ���"  ����#[  ����#[  ���"  �      !    ,��" 	U��" 
1��#[ 
1��#[ 	U��" 	U      !    ,��" +��" ��#[ ��#[ +��" +      !    ,��" ��" ���#[ ���#[ ��"       !    ,��" ���" x��#[ x��#[ ���" �      !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��2� ��2� ���3� ���3� ��2�       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��<� ��<� ���=� ���=� ��<�       !    ,��+� ���+� x��,� x��,� ���+� �      !    ,��%� +��%� ��&� ��&� +��%� +      !    ,��) +��) ��)� ��)� +��) +      !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��0� ���0� x��1k x��1k ���0� �      !    ,��%� 	U��%� 
1��&� 
1��&� 	U��%� 	U      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��5? ���5? x��6 x��6 ���5? �      !    ,��>� ���>� x��?{ x��?{ ���>� �      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��%� 	U��%� 
1��&� 
1��&� 	U��%� 	U      !    ,��0� ���0� x��1k x��1k ���0� �      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��) +��) ��)� ��)� +��) +      !    ,��%� +��%� ��&� ��&� +��%� +      !    ,��+� ���+� x��,� x��,� ���+� �      !    ,��<� ��<� ���=� ���=� ��<�       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��2� ��2� ���3� ���3� ��2�       !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��) ��) ���)� ���)� ��)       !    ,��%� ��%� ���&� ���&� ��%�       !    ,��'/ ���'/ x��( x��( ���'/ �      !    ,��9� ���9� x��:� x��:� ���9� �      !    ,��9� ���9� x��:� x��:� ���9� �      !    ,��'/ ���'/ x��( x��( ���'/ �      !    ,��%� ��%� ���&� ���&� ��%�       !    ,��) ��) ���)� ���)� ��)       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��>� ���>� x��?{ x��?{ ���>� �      !    ,��5? ���5? x��6 x��6 ���5? �      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��7 ��7 ���  ���  ��7       !    ,��� ���� x��� x��� ���� �      !    ,��o ���o x��K x��K ���o �      !    ,�� ��� x��� x��� ��� �      !    ,��� ���� x��� x��� ���� �      !    ,�� ��� x��� x��� ��� �      !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��_ 	U��_ 
1��; 
1��; 	U��_ 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��? ��? ���	 ���	 ��?       !    ,��� ��� ���c ���c ���       !    ,��� ��� ���� ���� ���       !    ,�� �� ���� ���� ��       !    ,��? +��? ��	 ��	 +��? +      !    ,��� +��� ��c ��c +��� +      !    ,��� +��� ��� ��� +��� +      !    ,�� +�� ��� ��� +�� +      !    ,��_ +��_ ��; ��; +��_ +      !    ,�� ��� x��� x��� ��� �      !    ,��� +��� ��� ��� +��� +      !    ,��_ ���_ x��; x��; ���_ �      !    ,��� +��� ��� ��� +��� +      !    ,��_ +��_ ��; ��; +��_ +      !    ,�� +�� ��� ��� +�� +      !    ,��� +��� ��� ��� +��� +      !    ,��� +��� ��c ��c +��� +      !    ,��? +��? ��	 ��	 +��? +      !    ,�� �� ���� ���� ��       !    ,��� ��� ���� ���� ���       !    ,��� ��� ���c ���c ���       !    ,��? ��? ���	 ���	 ��?       !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��_ 	U��_ 
1��; 
1��; 	U��_ 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,�� ��� x��� x��� ��� �      !    ,��� ���� x��� x��� ���� �      !    ,�� ��� x��� x��� ��� �      !    ,��o ���o x��K x��K ���o �      !    ,��� ���� x��� x��� ���� �      !    ,��7 ��7 ���  ���  ��7       !    ,��� ��� ���� ���� ���       !    ,��� ��� ���� ���� ���       !    ,��_ ��_ ���; ���; ��_       !    ,��7 +��7 ��  ��  +��7 +      !    ,��� +��� ��� ��� +��� +      !    ,��_ ���_ x��; x��; ���_ �      !    ,��� +��� ��� ��� +��� +      !    ,�� ��� x��� x��� ��� �      !    ,��7 +��7 ��  ��  +��7 +      !    ,��_ ��_ ���; ���; ��_       !    ,��� ��� ���� ���� ���       !    ,��� ��� ���� ���� ���       !    ,��  ���  �����  �����  ���  �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��� ���� ���� ���� ���� �      !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��W ���W ���3 ���3 ���W �      !    ,��� ���� ���{ ���{ ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��K ���K ���' ���' ���K �      !    ,��� ���� ���o ���o ���� �      !    ,�� � ��� � ���!� ���!� ��� � �      !    ,��  ���  �����  �����  ���  �      !    ,���  ����  �����  �����  ����  �      !    ,��o  ���o  ����K  ����K  ���o  �      !    ,�� ��� ���� ���� ��� �      !    ,��� ���� ���� ���� ���� �      !    ,��� ���� ���� ���� ���� �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��  ���  �����  �����  ���  �      !    ,��	� ���	� ���
� ���
� ���	� �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,��o  ���o  ����K  ����K  ���o  �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,�� � ��� � ���!� ���!� ��� � �      !    ,��� ���� ���o ���o ���� �      !    ,��K ���K ���' ���' ���K �      !    ,�� ��� ���� ���� ��� �      !    ,��� ���� ���{ ���{ ���� �      !    ,��W ���W ���3 ���3 ���W �      !    ,��  ���  �����  �����  ���  �      !    ,���  ����  �����  �����  ����  �      !    ,��	� ���	� ���
� ���
� ���	� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��3_ ���3_ ���4; ���4; ���3_ �      !    ,��9�  ���9�  ����:�  ����:�  ���9�  �      !    ,��5?  ���5?  ����6  ����6  ���5?  �      !    ,��0�  ���0�  ����1k  ����1k  ���0�  �      !    ,��+�  ���+�  ����,�  ����,�  ���+�  �      !    ,��'/  ���'/  ����(  ����(  ���'/  �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��'k ���'k ���(G ���(G ���'k �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��9� ���9� ���:� ���:� ���9� �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��-. ���-. ���.
 ���.
 ���-. �      !    ,��;W ���;W ���<3 ���<3 ���;W �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��'k ���'k ���(G ���(G ���'k �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��'/  ���'/  ����(  ����(  ���'/  �      !    ,��+�  ���+�  ����,�  ����,�  ���+�  �      !    ,��0�  ���0�  ����1k  ����1k  ���0�  �      !    ,��5?  ���5?  ����6  ����6  ���5?  �      !    ,��9�  ���9�  ����:�  ����:�  ���9�  �      !    ,��3_ ���3_ ���4; ���4; ���3_ �      !    ,��;W ���;W ���<3 ���<3 ���;W �      !    ,��-. ���-. ���.
 ���.
 ���-. �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��9� ���9� ���:� ���:� ���9� �      "    ,�� ��� G��! G��! ��� �      "    ,��K ���K ���O ���O ���K �      "    ,��"k ���"k /��#o /��#o ���"k �      "    ,��� ���� ���&� ���&� ���� �      "    ,�� � ��� � ���+� ���+� ��� � �      "    ,��2  �K��2  O��%  O��%  �K��2  �K      "    ,��/� ���/� ���0� ���0� ���/� �      "    ,��=� ���=� G��>� G��>� ���=� �      "    ,���  �����  �[��A  �[��A  �����  ��      "    ,��=� ���=� G��>� G��>� ���=� �      "    ,��/� ���/� ���0� ���0� ���/� �      "    ,��2  �K��2  O��%  O��%  �K��2  �K      "    ,�� � ��� � ���+� ���+� ��� � �      "    ,��� ���� ���&� ���&� ���� �      "    ,��"k ���"k ���#o ���#o ���"k �      "    ,��K ���K ���O ���O ���K �      "    ,�� ��� G��! G��! ��� �      "    ,��� ���� m��A m��A ���� �      "    ,��6 ���6 ���7 ���7 ���6 �      "    ,��%� ���%� ���&� ���&� ���%� �      "    ,��%� ���%� ���&� ���&� ���%� �      "    ,��6 ���6 ���7 ���7 ���6 �      "    ,��� ���� ��� ��� ���� �      "    ,��� ���� ��� ��� ���� �      "    ,��� ���� ���� ���� ���� �      "    ,��� ���� ���� ���� ���� �      "    ,��,C G��,C /��-G /��-G G��,C G      "    ,��(o ���(o ���*� ���*� ���(o �      "    ,��9c G��9c /��:g /��:g G��9c G      "    ,��<� 	K��<� ���=� ���=� 	K��<� 	K      "    ,��2� G��2� /��3� /��3� G��2� G      "    ,��2� G��2� ���3� ���3� G��2� G      "    ,��9c G��9c ���:g ���:g G��9c G      "    ,��<� G��<� 	K��>� 	K��>� G��<� G      "    ,��<� 	K��<� ���=� ���=� 	K��<� 	K      "    ,��<� G��<� 	K��>� 	K��>� G��<� G      "    ,��(o ���(o ���*� ���*� ���(o �      "    ,��,C G��,C ���-G ���-G G��,C G      "    ,��� ���� ��� � ��� � ���� �      "    ,��� G��� /��� /��� G��� G      "    ,��� G��� ���� ���� G��� G      "    ,��& 	K��& ���	* ���	* 	K��& 	K      "    ,��s G��s /��w /��w G��s G      "    ,�� G�� /�� /�� G�� G      "    ,��� ���� ��� � ��� � ���� �      "    ,�� G�� ��� ��� G�� G      "    ,��s G��s ���w ���w G��s G      "    ,�� G�� 	K��	* 	K��	* G�� G      "    ,��& 	K��& ���	* ���	* 	K��& 	K      "    ,�� G�� 	K��	* 	K��	* G�� G      "    ,��> }��> ���� ���� }��> }      "    ,��> }��> ���� ���� }��> }      "    ,��2  O��2 ���6 ���6  O��2  O      "    ,��� E��� ���� ���� E��� E      "    ,��� ?��� y�� y�� ?��� ?      "    ,�� � ?�� � ���!� ���!� ?�� � ?      "    ,��
�  �[��
� ���� ����  �[��
�  �[      "    ,��>  ���> }��B }��B  ���>  �      "    ,��	C O��	C /��
� /��
� O��	C O      "    ,��( ���( ���! ���! ���( �      "    ,��� E��� ���� ���� E��� E      "    ,�� ��� ���� ���� ��� �      "    ,��>  ���> }��B }��B  ���>  �      "    ,��
�  �[��
� ���� ����  �[��
�  �[      "    ,���  ���� ���� ����  ����  �      "    ,�� ��� ���� ���� ��� �      "    ,���  ���� ���� ����  ����  �      "    ,��	C O��	C /��
� /��
� O��	C O      "    ,��( ���( ���! ���! ���( �      "    ,���  �[��� ���� ����  �[���  �[      "    ,�� � ?�� � ���!� ���!� ?�� � ?      "    ,��� ?��� y�� y�� ?��� ?      "    ,��2  O��2 ���6 ���6  O��2  O      "    ,��7  ���7 ��� ���  ���7  �      "    ,���  �[��� ���� ����  �[���  �[      "    ,��7  ���7 ��� ���  ���7  �      "    ,��6 E��6 ���7� ���7� E��6 E      "    ,��6 E��6 ���7� ���7� E��6 E      "    ,��=� ���=� ���?� ���?� ���=� �      "    ,��6�  ���6� E��7� E��7�  ���6�  �      "    ,��3K  �[��3K ���4O ���4O  �[��3K  �[      "    ,��-[  ���-[ ���0� ���0�  ���-[  �      "    ,��'R  �[��'R ���(V ���(V  �[��'R  �[      "    ,��:� O��:� H��<� H��<� O��:� O      "    ,��:� O��:� H��<� H��<� O��:� O      "    ,��*�  ���*� ���+� ���+�  ���*�  �      "    ,��-[  ���-[ ���0� ���0�  ���-[  �      "    ,��3K  �[��3K ���4O ���4O  �[��3K  �[      "    ,��6�  ���6� E��7� E��7�  ���6�  �      "    ,��=� ���=� ���?� ���?� ���=� �      "    ,��9�  �[��9� ���:� ���:�  �[��9�  �[      "    ,��*�  ���*� ���+� ���+�  ���*�  �      "    ,��'R  �[��'R ���(V ���(V  �[��'R  �[      "    ,��=# ���=# ���>� ���>� ���=# �      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��=#  ���=# ���>' ���>'  ���=#  �      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��,� E��,� ���.� ���.� E��,� E      "    ,��=#  ���=# ���>' ���>'  ���=#  �      "    ,��=# ���=# ���>� ���>� ���=# �      "    ,��,� E��,� ���.� ���.� E��,� E      "    ,��9�  �[��9� ���:� ���:�  �[��9�  �[      #    ,��# ��# �� ' �� ' ��#       #    ,��(� ��(� ��)� ��)� ��(�       #    ,��# 
��# �� ' �� ' 
��# 
      #    ,��(� 
��(� ��)� ��)� 
��(� 
      #    ,��� ���� ���� ���� ���� �      #    ,��	� ���	� ���
� ���
� ���	� �      #    ,��u ��u ��y ��y ��u       #    ,��� ���� ���� ���� ���� �      #    ,��- ���- ���. ���. ���- �      #    ,��6\ ��6\ ��7` ��7` ��6\       #    ,��;C ���;C ���<G ���<G ���;C �      #    ,��>; ���>; ���?? ���?? ���>; �      #    ,��� ���� ���� ���� ���� �      #    ,�� ��� ���� ���� ��� �      #    ,��/1 ���/1 ���05 ���05 ���/1 �      #    ,��/1 ���/1 ���05 ���05 ���/1 �      #    ,�� ��� ���� ���� ��� �      #    ,��� ���� ���� ���� ���� �      #    ,��>; ���>; ���?? ���?? ���>; �      #    ,��;C ���;C ���<G ���<G ���;C �      #    ,��6\ ��6\ ��7` ��7` ��6\       #    ,��- ���- ���. ���. ���- �      #    ,��� ���� ���� ���� ���� �      #    ,��u ��u ��y ��y ��u       #    ,��	� ���	� ���
� ���
� ���	� �      #    ,��� ���� ���� ���� ���� �      #    ,��(� 
��(� ��)� ��)� 
��(� 
      #    ,��# 
��# �� ' �� ' 
��# 
      #    ,��(� ��(� ��)� ��)� ��(�       #    ,��# ��# �� ' �� ' ��#       $    ,��k *��k ��� � ��� � *��k *      $    ,��(o *��(o ���*� ���*� *��(o *      $    ,��k 
���k *��*� *��*� 
���k 
�      $    ,��k ���k 
��� � 
��� � ���k �      $    ,��(o ���(o 
���*� 
���*� ���(o �      $    ,��	C /��	C ���
o ���
o /��	C /      $    ,��( ���( ��� ��� ���( �      $    ,��	C O��	C /��
� /��
� O��	C O      $    ,��> ���> ���� ���� ���> �      $    ,��� ���� ���O ���O ���� �      $    ,��> ���> ���O ���O ���> �      $    ,��	C ���	C O��
o O��
o ���	C �      $    ,��> }��> ���� ���� }��> }      $    ,��� E��� ���O ���O E��� E      $    ,��7 ���7 ��� ��� ���7 �      $    ,��k y��k ���� ���� y��k y      $    ,��,� q��,� ���.� ���.� q��,� q      $    ,��6 q��6 ���7� ���7� q��6 q      $    ,��;k H��;k ���<� ���<� H��;k H      $    ,��,� E��,� q��7� q��7� E��,� E      $    ,��:� O��:� H��<� H��<� O��:� O      $    ,��	C  ���	C ��� ���  ���	C  �      $    ,��� ?��� y�� y�� ?��� ?      $    ,��-[ ���-[ ���0� ���0� ���-[ �      $    ,��;k ���;k O��<� O��<� ���;k �      $    ,��=� ���=� ���?� ���?� ���=� �      $    ,��k  ���k ?��� ?���  ���k  �      $    ,��-[  ���-[ ���<� ���<�  ���-[  �      $    ,��-[  ���-[ ���<� ���<�  ���-[  �      $    ,��k  ���k ?��� ?���  ���k  �      $    ,��=� ���=� ���?� ���?� ���=� �      $    ,��;k ���;k O��<� O��<� ���;k �      $    ,��-[ ���-[ ���0� ���0� ���-[ �      $    ,��� ?��� y�� y�� ?��� ?      $    ,��	C  ���	C ��� ���  ���	C  �      $    ,��:� O��:� H��<� H��<� O��:� O      $    ,��,� E��,� q��7� q��7� E��,� E      $    ,��;k H��;k ���<� ���<� H��;k H      $    ,��6 q��6 ���7� ���7� q��6 q      $    ,��,� q��,� ���.� ���.� q��,� q      $    ,��k y��k ���� ���� y��k y      $    ,��7 ���7 ��� ��� ���7 �      $    ,��� E��� ���O ���O E��� E      $    ,��> }��> ���� ���� }��> }      $    ,��	C ���	C O��
o O��
o ���	C �      $    ,��> ���> ���O ���O ���> �      $    ,��� ���� ���O ���O ���� �      $    ,��> ���> ���� ���� ���> �      $    ,��	C O��	C /��
� /��
� O��	C O      $    ,��( ���( ��� ��� ���( �      $    ,��	C /��	C ���
o ���
o /��	C /      $    ,��(o ���(o 
���*� 
���*� ���(o �      $    ,��k ���k 
��� � 
��� � ���k �      $    ,��k 
���k *��*� *��*� 
���k 
�      $    ,��(o *��(o ���*� ���*� *��(o *      $    ,��k *��k ��� � ��� � *��k *      $  
      @Y������ ��� � L       $  
      @Y������ ��� J E       $  
      @Y������ ��? x G       "  
      @I�^5?|� ��7�  VDD       "  
      @I�^5?|� ��7�  �� VSS         
 ��� � A         
 ��B � B         
 ��B � B         
 ��� � A       