  X � 
    � 
     LIB  >A�7KƧ�9D�/��ZT � 
    � 
     gf180mcu_gp9t3v3__comp2_2         ,���� ����� m��K$ m��K$ ����� �          ,��!v ��!v ���$d ���$d ��!v           ,��!v  ����!v  �u��$d  �u��$d  ����!v  ��          ,��!v  ����!v  �u��$d  �u��$d  ����!v  ��          ,��!v ��!v ���$d ���$d ��!v           ,��!� G��!� ���-� ���-� G��!� G          ,��8� ��8� ���;� ���;� ��8�           ,��&& ��&& ���) ���) ��&&           ,��=� ��=� ���@� ���@� ��=�           ,��=� ��=� ���@� ���@� ��=�           ,��*� ��*� ���-� ���-� ��*�           ,��BF ��BF ���E4 ���E4 ��BF           ,��BF ��BF ���E4 ���E4 ��BF           ,��8� ��8� ���;� ���;� ��8�           ,��46 ��46 ���7$ ���7$ ��46           ,��/� ��/� ���2t ���2t ��/�           ,��*� ��*� ���-� ���-� ��*�           ,��&& ��&& ���) ���) ��&&           ,��/� ��/� ���2t ���2t ��/�           ,��8� G��8� ���D� ���D� G��8� G          ,��.� G��.� ���7� ���7� G��.� G          ,��46 ��46 ���7$ ���7$ ��46           ,��BF ��BF ���E4 ���E4 ��BF           ,��BF ��BF ���E4 ���E4 ��BF           ,��F� ��F� ���I� ���I� ��F�           ,��F� ��F� ���I� ���I� ��F�           ,��F� ��F� ���I� ���I� ��F�           ,��F� ��F� ���I� ���I� ��F�           ,��
 ��
 ���� ���� ��
           ,��
 ��
 ���� ���� ��
           ,��� ��� ���� ���� ���           ,�� �� ��� ��� ��           ,��f ��f ���T ���T ��f           ,��� ��� ���� ���� ���           ,��
 ��
 ���� ���� ��
           ,�� � �� � ���� ���� �� �           ,��V ��V ���D ���D ��V           ,��� ��� ���� ���� ���           ,��
 ��
 ���� ���� ��
           ,�� G�� ��� ��� G�� G          ,��/ G��/ ��� � ��� � G��/ G          ,��� ��� ���� ���� ���           ,��V ��V ���D ���D ��V           ,��f ��f ���T ���T ��f           ,�� � �� � ���� ���� �� �           ,���� ���� ����� ����� ����           ,���� ���� ����� ����� ����           ,��f  ����f  �u��T  �u��T  ����f  ��          ,���  �����  �u���  �u���  �����  ��          ,��V  ����V  �u��D  �u��D  ����V  ��          ,��V  ����V  �u��D  �u��D  ����V  ��          ,��
  ����
  �u���  �u���  ����
  ��          ,�� �  ��� � ���� ����  ��� �  �          ,���  �����  �u���  �u���  �����  ��          ,��  ����  �u��  �u��  ����  ��          ,��f  ����f  �u��T  �u��T  ����f  ��          ,���  �����  �u���  �u���  �����  ��          ,��
  ����
  �u���  �u���  ����
  ��          ,��
  ����
  �u���  �u���  ����
  ��          ,��V  ����V  �u��D  �u��D  ����V  ��          ,��V  ����V  �u��D  �u��D  ����V  ��          ,���  ���� ���7 ���7  ����  �          ,��c  ���c ���"W ���"W  ���c  �          ,��
  ����
  �u���  �u���  ����
  ��          ,���  �����  �u���  �u���  �����  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,��/�  ����/�  �u��2t  �u��2t  ����/�  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��BF  ����BF  �u��E4  �u��E4  ����BF  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��9O  ���9O ���EC ���EC  ���9O  �          ,��0�  ���0� ���8# ���8#  ���0�  �          ,��#�  ���#� ���/w ���/w  ���#�  �          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��46  ����46  �u��7$  �u��7$  ����46  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��46  ����46  �u��7$  �u��7$  ����46  ��          ,��/�  ����/�  �u��2t  �u��2t  ����/�  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��          ,��&&  ����&&  �u��)  �u��)  ����&&  ��          ,��&&  ����&&  �u��)  �u��)  ����&&  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��           4���V k���V '���V m��J� m��J� k���V k           ,�� ��� ���U ���U ��� �           ,��� ���� ��� ��� ���� �           ,��� ���� ���!! ���!! ���� �           ,��  ����  ����U  ����U  ����  ��           ,���  �����  ����  ����  �����  ��           ,���  �����  ����!!  ����!!  �����  ��           ,���  �����  ����!!  ����!!  �����  ��           ,���  �����  ����  ����  �����  ��           ,��  ����  ����U  ����U  ����  ��           ,��� ���� ���!! ���!! ���� �           ,��� ���� ��� ��� ���� �           ,�� ��� ���U ���U ��� �           ,��$� ���$� ���.A ���.A ���$� �           ,��1� ���1� ���6� ���6� ���1� �           ,��:� ���:� ���@� ���@� ���:� �           ,��$�  ����$�  ����.A  ����.A  ����$�  ��           ,��1�  ����1�  ����6�  ����6�  ����1�  ��           ,��:�  ����:�  ����@�  ����@�  ����:�  ��           ,��:�  ����:�  ����@�  ����@�  ����:�  ��           ,��1�  ����1�  ����6�  ����6�  ����1�  ��           ,��$�  ����$�  ����.A  ����.A  ����$�  ��           ,����  ������ ���F) ���F)  ������  ��           ,��:� ���:� ���@� ���@� ���:� �           ,��1� ���1� ���6� ���6� ���1� �           ,��$� ���$� ���.A ���.A ���$� �          ,��R  ����R  ����h  ����h  ����R  ��          ,��B  ����B  ����X  ����X  ����B  ��          ,��	�  ����	�  ����  ����  ����	�  ��          ,��8�  ����8�  ����;�  ����;�  ����8�  ��          ,��4"  ����4"  ����78  ����78  ����4"  ��          ,��/r  ����/r  ����2�  ����2�  ����/r  ��          ,��*�  ����*�  ����-�  ����-�  ����*�  ��          ,��&  ����&  ����)(  ����)(  ����&  ��          ,��!b  ����!b  ����$x  ����$x  ����!b  ��          ,���  �����  �����  �����  �����  ��          ,��  ����  ����  ����  ����  ��          ,��=�  ����=�  ����@�  ����@�  ����=�  ��          ,���  �����  �����  �����  �����  ��          ,��B2  ����B2  ����EH  ����EH  ����B2  ��          ,�� ) a�� ) ���E� ���E� a�� ) a          ,��F�  ����F�  ����I�  ����I�  ����F�  ��          ,�� �  ���� �  �����  �����  ���� �  ��          ,����  ������  ������  ������  ������  ��          ,��K ���K ���< ���< ���K �          ,��s ���s ���� ���� ���s �          ,��	� ��	� ���
� ���
� ��	�           ,��>� U��>� ��C' ��C' U��>� U          ,��6 '��6 ��7� ��7� '��6 '          ,��	C U��	C ��
� ��
� U��	C U          ,��� ���� ���� ���� ���� �          ,��# ��# ���O ���O ��#           ,��O ��O ��� ; ��� ; ��O           ,���  ����� }�� }��  �����  ��          ,��� }��� E��� E��� }��� }          ,��� U��� �� �� U��� U          ,���  ����� U��� U���  �����  ��          ,��(� U��(� ��3� ��3� U��(� U          ,��%' ��%' ���(o ���(o ��%'           ,��:� E��:� ���< ���< E��:� E          ,��A�  ����A� U��C' U��C'  ����A�  ��          ,��>; ��>; ���B� ���B� ��>;           ,��	C  ����	C  ����6  ����6  ����	C  ��          ,��A� ���A� ���B� ���B� ���A� �          ,��	C  ����	C  ����6  ����6  ����	C  ��          ,��:� E��:� ���< ���< E��:� E          ,��4�  ����4� ��6 ��6  ����4�  ��          ,��%�  ����%� U��&� U��&�  ����%�  ��          ,��#� U��#� ��&� ��&� U��#� U          ,��#� ��#� ���%' ���%' ��#�           ,��  ���� �� ; �� ;  ����  ��          ,��  ���� }��� }���  ����  ��          ,���  ����� }�� }��  �����  ��          ,��� E��� ��� ��� E��� E          ,��k ���k ���� ���� ���k �          ,��� ���� ��� ��� ���� �          ,��� ���� ���� ���� ���� �          ,���  ����� '��� '���  �����  ��          ,��	C  ����	C U��
o U��
o  ����	C  ��          ,��� ��� ���w ���w ���           ,��K ���K ���w ���w ���K �          ,���  ����� U��' U��'  �����  ��          ,��� ��� ��� ��� ���           ,��s ���s ���� ���� ���s �          ,��K ���K ���< ���< ���K �          ,��+ ��+ ���� ���� ��+           ,��+ ���+ ���W ���W ���+ �          ,���  ����� U��� U���  �����  ��          ,��� U��� ��' ��' U��� U          ,��(�  ����(� U��* U��*  ����(�  ��          ,��>; ���>; ���?g ���?g ���>; �          ,��>; ��>; ��?� ��?� ��>;           ,��:� }��:� E��<� E��<� }��:� }          ,��;k  ����;k }��<� }��<�  ����;k  ��          ,��>�  ����>� U��?� U��?�  ����>�  ��          ,��;k  ����;k }��<� }��<�  ����;k  ��          ,��:� }��:� E��<� E��<� }��:� }          ,��2�  ����2� U��3� U��3�  ����2�  ��          ,��,/  ����,/ U��-[ U��-[  ����,/  ��          ,��/� ��/� ��1� ��1� ��/�           ,��4c ��4c ���6 ���6 ��4c           ,��4c ���4c ���5� ���5� ���4c �          ,��*� ��*� ���2G ���2G ��*�           ,��1 ���1 ���2G ���2G ���1 �          ,��*� ���*� ���+� ���+� ���*� �          ,��'C ���'C ���(o ���(o ���'C �          ,�� '�� ��� ��� '�� '      !    ,��" ~��" Z��#[ Z��#[ ~��" ~      !    ,��"  �&��"  ���#[  ���#[  �&��"  �&      !    ,��"  �&��"  ���#[  ���#[  �&��"  �&      !    ,��" 	U��" 
1��#[ 
1��#[ 	U��" 	U      !    ,��" +��" ��#[ ��#[ +��" +      !    ,��" ��" ���#[ ���#[ ��"       !    ,��" ~��" Z��#[ Z��#[ ~��" ~      !    ,��%� ��%� ���&� ���&� ��%�       !    ,��%� +��%� ��&� ��&� +��%� +      !    ,��%� 	U��%� 
1��&� 
1��&� 	U��%� 	U      !    ,��+� ~��+� Z��,� Z��,� ~��+� ~      !    ,��) +��) ��)� ��)� +��) +      !    ,��0� ~��0� Z��1k Z��1k ~��0� ~      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��5? ~��5? Z��6 Z��6 ~��5? ~      !    ,��>� ~��>� Z��?{ Z��?{ ~��>� ~      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��0� ~��0� Z��1k Z��1k ~��0� ~      !    ,��) +��) ��)� ��)� +��) +      !    ,��+� ~��+� Z��,� Z��,� ~��+� ~      !    ,��) ��) ���)� ���)� ��)       !    ,��'/ ~��'/ Z��( Z��( ~��'/ ~      !    ,��9� ~��9� Z��:� Z��:� ~��9� ~      !    ,��9� ~��9� Z��:� Z��:� ~��9� ~      !    ,��'/ ~��'/ Z��( Z��( ~��'/ ~      !    ,��) ��) ���)� ���)� ��)       !    ,��>� ~��>� Z��?{ Z��?{ ~��>� ~      !    ,��5? ~��5? Z��6 Z��6 ~��5? ~      !    ,��CO ~��CO Z��D+ Z��D+ ~��CO ~      !    ,��CO ~��CO Z��D+ Z��D+ ~��CO ~      !    ,��CO ~��CO Z��D+ Z��D+ ~��CO ~      !    ,��CO ~��CO Z��D+ Z��D+ ~��CO ~      !    ,��G� ~��G� Z��H� Z��H� ~��G� ~      !    ,��G� ~��G� Z��H� Z��H� ~��G� ~      !    ,��G� ~��G� Z��H� Z��H� ~��G� ~      !    ,��G� ~��G� Z��H� Z��H� ~��G� ~      !    ,��CO 	U��CO 
1��D+ 
1��D+ 	U��CO 	U      !    ,��CO ��CO ���D+ ���D+ ��CO       !    ,��CO +��CO ��D+ ��D+ +��CO +      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��@ 	U��@ 
1��@� 
1��@� 	U��@ 	U      !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��2� ��2� ���3� ���3� ��2�       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��<� ��<� ���=� ���=� ��<�       !    ,��@ ��@ ���@� ���@� ��@       !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��@ +��@ ��@� ��@� +��@ +      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��@ 	U��@ 
1��@� 
1��@� 	U��@ 	U      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��@ +��@ ��@� ��@� +��@ +      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��@ ��@ ���@� ���@� ��@       !    ,��<� ��<� ���=� ���=� ��<�       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��2� ��2� ���3� ���3� ��2�       !    ,�� ~�� Z��� Z��� ~�� ~      !    ,��7 +��7 ��  ��  +��7 +      !    ,�� �� ���� ���� ��       !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� ��� ���� ���� ���       !    ,��7 ��7 ���  ���  ��7       !    ,��� ~��� Z��� Z��� ~��� ~      !    ,��o ~��o Z��K Z��K ~��o ~      !    ,�� ~�� Z��� Z��� ~�� ~      !    ,��� ~��� Z��� Z��� ~��� ~      !    ,��� +��� ��� ��� +��� +      !    ,��� ��� ���� ���� ���       !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��� ~��� Z��� Z��� ~��� ~      !    ,��� ~��� Z��� Z��� ~��� ~      !    ,���� ~���� Z���� Z���� ~���� ~      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��� ��� ���� ���� ���       !    ,��? ��? ���	 ���	 ��?       !    ,��� ��� ���c ���c ���       !    ,��� ��� ���� ���� ���       !    ,��� +��� ��� ��� +��� +      !    ,��? +��? ��	 ��	 +��? +      !    ,��� +��� ��c ��c +��� +      !    ,��� +��� ��� ��� +��� +      !    ,�� +�� ��� ��� +�� +      !    ,�� ~�� Z��� Z��� ~�� ~      !    ,��� +��� ��� ��� +��� +      !    ,��_ ~��_ Z��; Z��; ~��_ ~      !    ,�� ~�� Z��� Z��� ~�� ~      !    ,�� +�� ��� ��� +�� +      !    ,��_ +��_ ��; ��; +��_ +      !    ,��� +��� ��c ��c +��� +      !    ,��? +��? ��	 ��	 +��? +      !    ,��� +��� ��� ��� +��� +      !    ,��_ ��_ ���; ���; ��_       !    ,��� ��� ���c ���c ���       !    ,��? ��? ���	 ���	 ��?       !    ,��� ��� ���� ���� ���       !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��_ 	U��_ 
1��; 
1��; 	U��_ 	U      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� ~�� Z��� Z��� ~�� ~      !    ,��� ~��� Z��� Z��� ~��� ~      !    ,�� ~�� Z��� Z��� ~�� ~      !    ,��o ~��o Z��K Z��K ~��o ~      !    ,��� ~��� Z��� Z��� ~��� ~      !    ,��7 ��7 ���  ���  ��7       !    ,��� ��� ���� ���� ���       !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,�� �� ���� ���� ��       !    ,��7 +��7 ��  ��  +��7 +      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��_ ~��_ Z��; Z��; ~��_ ~      !    ,��� +��� ��� ��� +��� +      !    ,���� ~���� Z���� Z���� ~���� ~      !    ,���  �&���  ����  ����  �&���  �&      !    ,��  �&��  ����  ����  �&��  �&      !    ,��� ���� ���o ���o ���� �      !    ,��K ���K ���' ���' ���K �      !    ,�� � ��� � ���!� ���!� ��� � �      !    ,��� ���� ���� ���� ���� �      !    ,��W ���W ���3 ���3 ���W �      !    ,�� ��� ���� ���� ��� �      !    ,��  �&��  ����  ����  �&��  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,��_ ���_ ���; ���; ���_ �      !    ,��  �&��  ����  ����  �&��  �&      !    ,��_  �&��_  ���;  ���;  �&��_  �&      !    ,��_  �&��_  ���;  ���;  �&��_  �&      !    ,�� ��� ���[ ���[ ��� �      !    ,��� ���� ���� ���� ���� �      !    ,��  �&��  ����  ����  �&��  �&      !    ,�� ��� ���� ���� ��� �      !    ,��W ���W ���3 ���3 ���W �      !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��7 ���7 ��� ��� ���7 �      !    ,���  �&���  ����  ����  �&���  �&      !    ,��o  �&��o  ���K  ���K  �&��o  �&      !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���[ ���[ ��� �      !    ,��_  �&��_  ���;  ���;  �&��_  �&      !    ,��� ���� ���o ���o ���� �      !    ,��_  �&��_  ���;  ���;  �&��_  �&      !    ,��  �&��  ����  ����  �&��  �&      !    ,��_ ���_ ���; ���; ���_ �      !    ,���  �&���  ����  ����  �&���  �&      !    ,��  �&��  ����  ����  �&��  �&      !    ,��o  �&��o  ���K  ���K  �&��o  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,���  �&���  ����  ����  �&���  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,����  �&����  �����  �����  �&����  �&      !    ,��_ ���_ ���; ���; ���_ �      !    ,��� ���� ���n ���n ���� �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��1C ���1C ���2 ���2 ���1C �      !    ,��C� ���C� ���D� ���D� ���C� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��9� ���9� ���:� ���:� ���9� �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��@ ���@ ���A[ ���A[ ���@ �      !    ,��0v ���0v ���1R ���1R ���0v �      !    ,��>� ���>� ���?{ ���?{ ���>� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��1C ���1C ���2 ���2 ���1C �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��>� ���>� ���?{ ���?{ ���>� �      !    ,��0v ���0v ���1R ���1R ���0v �      !    ,��@ ���@ ���A[ ���A[ ���@ �      !    ,��'k ���'k ���(G ���(G ���'k �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��CO  �&��CO  ���D+  ���D+  �&��CO  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��G�  �&��G�  ���H�  ���H�  �&��G�  �&      !    ,��>�  �&��>�  ���?{  ���?{  �&��>�  �&      !    ,��>�  �&��>�  ���?{  ���?{  �&��>�  �&      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��'/  �&��'/  ���(  ���(  �&��'/  �&      !    ,��+�  �&��+�  ���,�  ���,�  �&��+�  �&      !    ,��0�  �&��0�  ���1k  ���1k  �&��0�  �&      !    ,��5?  �&��5?  ���6  ���6  �&��5?  �&      !    ,��9�  �&��9�  ���:�  ���:�  �&��9�  �&      !    ,��>�  �&��>�  ���?{  ���?{  �&��>�  �&      !    ,��>�  �&��>�  ���?{  ���?{  �&��>�  �&      !    ,��9�  �&��9�  ���:�  ���:�  �&��9�  �&      !    ,��5?  �&��5?  ���6  ���6  �&��5?  �&      !    ,��0�  �&��0�  ���1k  ���1k  �&��0�  �&      !    ,��+�  �&��+�  ���,�  ���,�  �&��+�  �&      !    ,��'/  �&��'/  ���(  ���(  �&��'/  �&      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��9� ���9� ���:� ���:� ���9� �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��6� ���6� ���7j ���7j ���6� �      "    ,��� ���� G��� G��� ���� �      "    ,�� ��� ��� ��� ��� �      "    ,��%� ���%� ���&� ���&� ���%� �      "    ,��� ���� ���)� ���)� ���� �      "    ,��� :��� V��� V��� :��� :      "    ,����  ������  �[��K$  �[��K$  ������  ��      "    ,���  �K���  O��%  O��%  �K���  �K      "    ,��� ���� ���)� ���)� ���� �      "    ,��# ���# ��� ' ��� ' ���# �      "    ,�� ��� ��� ��� ��� �      "    ,��� /��� G��� G��� /��� /      "    ,���� ����� m��K$ m��K$ ����� �      "    ,��(� ���(� ���)� ���)� ���(� �      "    ,��(� ���(� ���)� ���)� ���(� �      "    ,��� E��� ���� ���� E��� E      "    ,��� ���� ��� ��� ���� �      "    ,��n ���n ���r ���r ���n �      "    ,��n ���n ���r ���r ���n �      "    ,��/� G��/� /��0� /��0� G��/� G      "    ,��C; G��C; ���D? ���D? G��C; G      "    ,��6 ���6 ���7 ���7 ���6 �      "    ,��<� G��<� ���=� ���=� G��<� G      "    ,��/� G��/� ���0� ���0� G��/� G      "    ,��"k ���"k ���#o ���#o ���"k �      "    ,�� ; :�� ; V��"W V��"W :�� ; :      "    ,��� 	K��� ���� ���� 	K��� 	K      "    ,��� G��� ���� ���� G��� G      "    ,��� ���� ���� ���� ���� �      "    ,��O ���O ���k ���k ���O �      "    ,��K G��K ���O ���O G��K G      "    ,��+ G��+ ���	/ ���	/ G��+ G      "    ,��� G��� 	K��� 	K��� G��� G      "    ,��� 	K��� ���� ���� 	K��� 	K      "    ,��� G��� 	K��� 	K��� G��� G      "    ,��
� }��
� ���r ���r }��
� }      "    ,��
� }��
� ���r ���r }��
� }      "    ,���  �[��� ���� ����  �[���  �[      "    ,��
�  ���
� }��� }���  ���
�  �      "    ,��� O��� /��� /��� O��� O      "    ,��� ���� O��� O��� ���� �      "    ,���  �[��� ���� ����  �[���  �[      "    ,��
�  ���
� }��� }���  ���
�  �      "    ,��k  ���k ���o ���o  ���k  �      "    ,��� ���� ���o ���o ���� �      "    ,��k  ���k ���o ���o  ���k  �      "    ,��� O��� /��� /��� O��� O      "    ,��� O��� /��� /��� O��� O      "    ,��C  �[��C ���G ���G  �[��C  �[      "    ,�� ?�� ���� ���� ?�� ?      "    ,���  O��� ���� ����  O���  O      "    ,���  ���� ���7 ���7  ����  �      "    ,��'W  �[��'W ���([ ���([  �[��'W  �[      "    ,���  ���� ���7 ���7  ����  �      "    ,��#  �[��# ���' ���'  �[��#  �[      "    ,��6�  �[��6� ���7� ���7�  �[��6�  �[      "    ,��-�  �[��-� ���.� ���.�  �[��-�  �[      "    ,��=#  �[��=# ���>' ���>'  �[��=#  �[      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��=#  �[��=# ���>' ���>'  �[��=#  �[      "    ,��C�  �[��C� ���D� ���D�  �[��C�  �[      "    ,��6 '��6 ���7� ���7� '��6 '      "    ,��@k ���@k ���A� ���A� ���@k �      "    ,��@k  ���@k ���Ao ���Ao  ���@k  �      "    ,��/� E��/� ���1� ���1� E��/� E      "    ,��@k  ���@k ���Ao ���Ao  ���@k  �      "    ,��@k ���@k ���A� ���A� ���@k �      "    ,��@� ���@� O��A� O��A� ���@� �      "    ,��9�  ���9� E��:� E��:�  ���9�  �      "    ,��0�  ���0� ���3� ���3�  ���0�  �      "    ,��*�  ���*� ���+� ���+�  ���*�  �      "    ,��>; O��>; H��?� H��?� O��>; O      "    ,��>; O��>; H��?� H��?� O��>; O      "    ,��0�  ���0� ���3� ���3�  ���0�  �      "    ,��9�  ���9� E��:� E��:�  ���9�  �      "    ,��@� O��@� H��B� H��B� O��@� O      "    ,��9c E��9c ���:� ���:� E��9c E      "    ,��9c E��9c ���:� ���:� E��9c E      "    ,��+� ���+� ���-� ���-� ���+� �      "    ,��?� G��?� 	K��A� 	K��A� G��?� G      "    ,��?� 	K��?� ���@� ���@� 	K��?� 	K      "    ,��?� G��?� 	K��A� 	K��A� G��?� G      "    ,��?� 	K��?� ���@� ���@� 	K��?� 	K      "    ,��+� ���+� ���-� ���-� ���+� �      "    ,��9c ���9c ���:g ���:g ���9c �      "    ,��9c ���9c ���:g ���:g ���9c �      "    ,��2� ���2� ���3� ���3� ���2� �      "    ,��@� H��@� G��A� G��A� H��@� H      "    ,��2� ���2� ���3� ���3� ���2� �      "    ,�� ��� ���+� ���+� ��� �      "    ,�� '�� ���� ���� '�� '      #    ,��� ��� ��� ��� ���       #    ,��� 
��� ��� ��� 
��� 
      #    ,��K ���K ���O ���O ���K �      #    ,��- ��- ��1 ��1 ��-       #    ,�� � ��� � ���!� ���!� ��� � �      #    ,��� ��� ��� ��� ���       #    ,��K ���K ���O ���O ���K �      #    ,��7 ���7 ���; ���; ���7 �      #    ,��- ��- ��1 ��1 ��-       #    ,��K ���K ���O ���O ���K �      #    ,��X ���X ���\ ���\ ���X �      #    ,��,C ��,C ��-G ��-G ��,C       #    ,��,C 
��,C ��-G ��-G 
��,C 
      #    ,��0b ���0b ���1f ���1f ���0b �      #    ,��9� ��9� ��:� ��:� ��9�       #    ,��>� ���>� ���?� ���?� ���>� �      #    ,��A� ���A� ���B� ���B� ���A� �      #    ,��1/ &��1/ *��23 *��23 &��1/ &      #    ,��A� ���A� ���B� ���B� ���A� �      #    ,��>� ���>� ���?� ���?� ���>� �      #    ,��9� ��9� ��:� ��:� ��9�       #    ,��0b ���0b ���1f ���1f ���0b �      #    ,��,C 
��,C ��-G ��-G 
��,C 
      #    ,��,C ��,C ��-G ��-G ��,C       #    ,��X ���X ���\ ���\ ���X �      #    ,��[ ]��[ a��_ a��_ ]��[ ]      #    ,��6W ]��6W a��7[ a��7[ ]��6W ]   	   $    !    , $��1H ���1H K��9� K��9� �   	   $    !    , $��� I��� K��U K��U X      $    ,��� E��� ���� ���� E��� E      $    ,��/� E��/� ��1� ��1� E��/� E      $    ,��� O��� /��� /��� O��� O      $    ,��
� ���
� ���r ���r ���
� �      $    ,��� :��� V��� V��� :��� :      $    ,�� ; :�� ; V��"W V��"W :�� ; :      $    ,��� ���� O��' O��' ���� �      $    ,��6 ��6 ���7� ���7� ��6       $    ,��� :��� V��"W V��"W :��� :      $    ,�� �� ���� ���� ��       $    ,���  �����  ���7  ���7  �����  ��      $    ,��  ��� ���7 ���7  ���  �      $    ,���  ���� O��' O��'  ����  �      $    ,��
� I��
� ���r ���r I��
� I      $    ,��� O��� /��� /��� O��� O      $    ,��� O��� /��� /��� O��� O      $    ,��� /��� ���� ���� /��� /      $    ,��O V��O 
���k 
���k V��O V      $    ,��O *��O ���k ���k *��O *      $    ,��+� *��+� ���-� ���-� *��+� *      $    ,��+� ���+� 
���-� 
���-� ���+� �      $    ,��>� H��>� ���?� ���?� H��>� H      $    ,��>; O��>; H��?� H��?� O��>; O      $    ,��>� ���>� O��?� O��?� ���>� �      $    ,��0�  ���0� ���?� ���?�  ���0�  �      $    ,��0�  ���0� ���?� ���?�  ���0�  �      $    ,��@� O��@� H��B� H��B� O��@� O      $    ,��>� ���>� O��?� O��?� ���>� �      $    ,��0� ���0� ���3� ���3� ���0� �      $    ,��>; O��>; H��?� H��?� O��>; O      $    ,��>� H��>� ���?� ���?� H��>� H      $    ,��9c E��9c ���:� ���:� E��9c E      $    ,��+� ���+� 
���-� 
���-� ���+� �      $    ,��O 
���O *��-� *��-� 
���O 
�      $    ,��+� *��+� ���-� ���-� *��+� *      $  
   ��  � B       $  
   ��6� 9 A       $  
      @Y������ ��AL | G       $  
      @Y������ ��� : L       $  
      @Y������ ��� J E       "  
      @I�^5?|� ��7�  VDD       "  
      @I�^5?|� ��7�  �� VSS       