magic
tech gf180mcuD
magscale 1 10
timestamp 1755786031
<< nwell >>
rect -1662 -417 1299 530
<< nmos >>
rect -1454 -782 -1394 -612
rect -1284 -782 -1224 -612
rect -1114 -782 -1054 -612
rect -790 -782 -730 -612
rect -470 -782 -410 -612
rect -300 -782 -240 -612
rect -130 -782 -70 -612
rect 40 -782 100 -612
rect 360 -782 420 -612
rect 684 -782 744 -612
rect 854 -782 914 -612
rect 1024 -782 1084 -612
<< pmos >>
rect -1454 -252 -1394 88
rect -1284 -252 -1224 88
rect -1114 -252 -1054 88
rect -790 -252 -730 88
rect -470 -252 -410 88
rect -300 -252 -240 88
rect -130 -252 -70 88
rect 40 -252 100 88
rect 360 -252 420 88
rect 684 -252 744 88
rect 854 -252 914 88
rect 1024 -252 1084 88
<< ndiff >>
rect -1554 -672 -1454 -612
rect -1554 -718 -1531 -672
rect -1485 -718 -1454 -672
rect -1554 -782 -1454 -718
rect -1394 -674 -1284 -612
rect -1394 -720 -1364 -674
rect -1318 -720 -1284 -674
rect -1394 -782 -1284 -720
rect -1224 -782 -1114 -612
rect -1054 -679 -954 -612
rect -1054 -725 -1023 -679
rect -977 -725 -954 -679
rect -1054 -782 -954 -725
rect -894 -677 -790 -612
rect -894 -723 -867 -677
rect -821 -723 -790 -677
rect -894 -782 -790 -723
rect -730 -677 -630 -612
rect -730 -723 -699 -677
rect -653 -723 -630 -677
rect -730 -782 -630 -723
rect -570 -677 -470 -612
rect -570 -723 -547 -677
rect -501 -723 -470 -677
rect -570 -782 -470 -723
rect -410 -680 -300 -612
rect -410 -726 -378 -680
rect -332 -726 -300 -680
rect -410 -782 -300 -726
rect -240 -782 -130 -612
rect -70 -677 40 -612
rect -70 -723 -38 -677
rect 8 -723 40 -677
rect -70 -782 40 -723
rect 100 -677 200 -612
rect 100 -723 131 -677
rect 177 -723 200 -677
rect 100 -782 200 -723
rect 260 -677 360 -612
rect 260 -723 283 -677
rect 329 -723 360 -677
rect 260 -782 360 -723
rect 420 -678 524 -612
rect 420 -724 451 -678
rect 497 -724 524 -678
rect 420 -782 524 -724
rect 584 -674 684 -612
rect 584 -720 608 -674
rect 654 -720 684 -674
rect 584 -782 684 -720
rect 744 -782 854 -612
rect 914 -673 1024 -612
rect 914 -719 946 -673
rect 992 -719 1024 -673
rect 914 -782 1024 -719
rect 1084 -677 1184 -612
rect 1084 -723 1115 -677
rect 1161 -723 1184 -677
rect 1084 -782 1184 -723
<< pdiff >>
rect -1554 46 -1454 88
rect -1554 -200 -1531 46
rect -1485 -200 -1454 46
rect -1554 -252 -1454 -200
rect -1394 46 -1284 88
rect -1394 -200 -1364 46
rect -1318 -200 -1284 46
rect -1394 -252 -1284 -200
rect -1224 46 -1114 88
rect -1224 -200 -1192 46
rect -1146 -200 -1114 46
rect -1224 -252 -1114 -200
rect -1054 46 -954 88
rect -1054 -200 -1023 46
rect -977 -200 -954 46
rect -1054 -252 -954 -200
rect -894 46 -790 88
rect -894 -200 -867 46
rect -821 -200 -790 46
rect -894 -252 -790 -200
rect -730 46 -470 88
rect -730 -200 -631 46
rect -585 -200 -470 46
rect -730 -252 -470 -200
rect -410 46 -300 88
rect -410 -200 -378 46
rect -332 -200 -300 46
rect -410 -252 -300 -200
rect -240 46 -130 88
rect -240 -200 -208 46
rect -162 -200 -130 46
rect -240 -252 -130 -200
rect -70 46 40 88
rect -70 -200 -38 46
rect 8 -200 40 46
rect -70 -252 40 -200
rect 100 46 360 88
rect 100 -200 205 46
rect 251 -200 360 46
rect 100 -252 360 -200
rect 420 46 524 88
rect 420 -200 451 46
rect 497 -200 524 46
rect 420 -252 524 -200
rect 584 46 684 88
rect 584 -200 608 46
rect 654 -200 684 46
rect 584 -252 684 -200
rect 744 46 854 88
rect 744 -200 776 46
rect 822 -200 854 46
rect 744 -252 854 -200
rect 914 46 1024 88
rect 914 -200 946 46
rect 992 -200 1024 46
rect 914 -252 1024 -200
rect 1084 46 1184 88
rect 1084 -200 1115 46
rect 1161 -200 1184 46
rect 1084 -252 1184 -200
<< ndiffc >>
rect -1531 -718 -1485 -672
rect -1364 -720 -1318 -674
rect -1023 -725 -977 -679
rect -867 -723 -821 -677
rect -699 -723 -653 -677
rect -547 -723 -501 -677
rect -378 -726 -332 -680
rect -38 -723 8 -677
rect 131 -723 177 -677
rect 283 -723 329 -677
rect 451 -724 497 -678
rect 608 -720 654 -674
rect 946 -719 992 -673
rect 1115 -723 1161 -677
<< pdiffc >>
rect -1531 -200 -1485 46
rect -1364 -200 -1318 46
rect -1192 -200 -1146 46
rect -1023 -200 -977 46
rect -867 -200 -821 46
rect -631 -200 -585 46
rect -378 -200 -332 46
rect -208 -200 -162 46
rect -38 -200 8 46
rect 205 -200 251 46
rect 451 -200 497 46
rect 608 -200 654 46
rect 776 -200 822 46
rect 946 -200 992 46
rect 1115 -200 1161 46
<< psubdiff >>
rect -1570 -1074 -1420 -1052
rect -1570 -1120 -1518 -1074
rect -1472 -1120 -1420 -1074
rect -1570 -1142 -1420 -1120
rect -1330 -1074 -1180 -1052
rect -1330 -1120 -1278 -1074
rect -1232 -1120 -1180 -1074
rect -1330 -1142 -1180 -1120
rect -1090 -1074 -940 -1052
rect -1090 -1120 -1038 -1074
rect -992 -1120 -940 -1074
rect -1090 -1142 -940 -1120
rect -850 -1074 -700 -1052
rect -850 -1120 -798 -1074
rect -752 -1120 -700 -1074
rect -850 -1142 -700 -1120
rect -610 -1074 -460 -1052
rect -610 -1120 -558 -1074
rect -512 -1120 -460 -1074
rect -610 -1142 -460 -1120
rect -370 -1074 -220 -1052
rect -370 -1120 -318 -1074
rect -272 -1120 -220 -1074
rect -370 -1142 -220 -1120
rect -130 -1074 20 -1052
rect -130 -1120 -78 -1074
rect -32 -1120 20 -1074
rect -130 -1142 20 -1120
rect 110 -1074 260 -1052
rect 110 -1120 162 -1074
rect 208 -1120 260 -1074
rect 110 -1142 260 -1120
rect 350 -1074 500 -1052
rect 350 -1120 402 -1074
rect 448 -1120 500 -1074
rect 350 -1142 500 -1120
rect 590 -1074 740 -1052
rect 590 -1120 642 -1074
rect 688 -1120 740 -1074
rect 590 -1142 740 -1120
rect 830 -1074 980 -1052
rect 830 -1120 882 -1074
rect 928 -1120 980 -1074
rect 830 -1142 980 -1120
rect 1070 -1074 1220 -1052
rect 1070 -1120 1122 -1074
rect 1168 -1120 1220 -1074
rect 1070 -1142 1220 -1120
<< nsubdiff >>
rect -1570 426 -1420 448
rect -1570 380 -1518 426
rect -1472 380 -1420 426
rect -1570 358 -1420 380
rect -1330 426 -1180 448
rect -1330 380 -1278 426
rect -1232 380 -1180 426
rect -1330 358 -1180 380
rect -1090 426 -940 448
rect -1090 380 -1038 426
rect -992 380 -940 426
rect -1090 358 -940 380
rect -850 426 -700 448
rect -850 380 -798 426
rect -752 380 -700 426
rect -850 358 -700 380
rect -610 426 -460 448
rect -610 380 -558 426
rect -512 380 -460 426
rect -610 358 -460 380
rect -370 426 -220 448
rect -370 380 -318 426
rect -272 380 -220 426
rect -370 358 -220 380
rect -130 426 20 448
rect -130 380 -78 426
rect -32 380 20 426
rect -130 358 20 380
rect 110 426 260 448
rect 110 380 162 426
rect 208 380 260 426
rect 110 358 260 380
rect 350 426 500 448
rect 350 380 402 426
rect 448 380 500 426
rect 350 358 500 380
rect 590 426 740 448
rect 590 380 642 426
rect 688 380 740 426
rect 590 358 740 380
rect 830 426 980 448
rect 830 380 882 426
rect 928 380 980 426
rect 830 358 980 380
rect 1070 426 1220 448
rect 1070 380 1122 426
rect 1168 380 1220 426
rect 1070 358 1220 380
<< psubdiffcont >>
rect -1518 -1120 -1472 -1074
rect -1278 -1120 -1232 -1074
rect -1038 -1120 -992 -1074
rect -798 -1120 -752 -1074
rect -558 -1120 -512 -1074
rect -318 -1120 -272 -1074
rect -78 -1120 -32 -1074
rect 162 -1120 208 -1074
rect 402 -1120 448 -1074
rect 642 -1120 688 -1074
rect 882 -1120 928 -1074
rect 1122 -1120 1168 -1074
<< nsubdiffcont >>
rect -1518 380 -1472 426
rect -1278 380 -1232 426
rect -1038 380 -992 426
rect -798 380 -752 426
rect -558 380 -512 426
rect -318 380 -272 426
rect -78 380 -32 426
rect 162 380 208 426
rect 402 380 448 426
rect 642 380 688 426
rect 882 380 928 426
rect 1122 380 1168 426
<< polysilicon >>
rect -1284 288 100 338
rect -1454 88 -1394 138
rect -1284 88 -1224 288
rect -1114 188 -410 238
rect -1114 88 -1054 188
rect -790 88 -730 138
rect -470 88 -410 188
rect 40 188 100 288
rect 40 138 420 188
rect -300 88 -240 138
rect -130 88 -70 138
rect 40 88 100 138
rect 360 88 420 138
rect 684 88 744 138
rect 854 88 914 138
rect 1024 88 1084 138
rect -1454 -482 -1394 -252
rect -1454 -509 -1332 -482
rect -1454 -555 -1405 -509
rect -1359 -555 -1332 -509
rect -1454 -582 -1332 -555
rect -1454 -612 -1394 -582
rect -1284 -612 -1224 -252
rect -1114 -333 -1054 -252
rect -1114 -359 -972 -333
rect -1114 -405 -1045 -359
rect -999 -405 -972 -359
rect -1114 -432 -972 -405
rect -1114 -612 -1054 -432
rect -790 -612 -730 -252
rect -470 -612 -410 -252
rect -300 -612 -240 -252
rect -130 -612 -70 -252
rect 40 -612 100 -252
rect 360 -612 420 -252
rect 684 -302 744 -252
rect 624 -329 744 -302
rect 624 -375 651 -329
rect 697 -375 744 -329
rect 624 -402 744 -375
rect 684 -612 744 -402
rect 854 -612 914 -252
rect 1024 -472 1084 -252
rect 964 -499 1084 -472
rect 964 -545 991 -499
rect 1037 -545 1084 -499
rect 964 -572 1084 -545
rect 1024 -612 1084 -572
rect -1454 -832 -1394 -782
rect -1284 -832 -1224 -782
rect -1114 -832 -1054 -782
rect -790 -882 -730 -782
rect -470 -832 -410 -782
rect -300 -882 -240 -782
rect -790 -932 -240 -882
rect -130 -882 -70 -782
rect 40 -832 100 -782
rect 360 -832 420 -782
rect 684 -882 744 -782
rect -130 -932 744 -882
rect -300 -982 -240 -932
rect 854 -982 914 -782
rect 1024 -832 1084 -782
rect -300 -1032 914 -982
<< polycontact >>
rect -1405 -555 -1359 -509
rect -1045 -405 -999 -359
rect 651 -375 697 -329
rect 991 -545 1037 -499
<< metal1 >>
rect -1599 426 1250 498
rect -1599 380 -1518 426
rect -1472 380 -1278 426
rect -1232 380 -1038 426
rect -992 380 -798 426
rect -752 380 -558 426
rect -512 380 -318 426
rect -272 380 -78 426
rect -32 380 162 426
rect 208 380 402 426
rect 448 380 642 426
rect 688 380 882 426
rect 928 380 1122 426
rect 1168 380 1250 426
rect -1599 358 1250 380
rect -1534 46 -1482 88
rect -1534 -200 -1531 46
rect -1485 -200 -1482 46
rect -1534 -672 -1482 -200
rect -1367 46 -1315 358
rect -1367 -200 -1364 46
rect -1318 -200 -1315 46
rect -1367 -252 -1315 -200
rect -1193 46 -1141 87
rect -1193 -200 -1192 46
rect -1146 -200 -1141 46
rect -1193 -504 -1141 -200
rect -1026 46 -974 358
rect -1026 -200 -1023 46
rect -977 -200 -974 46
rect -1026 -252 -974 -200
rect -870 46 -818 88
rect -870 -200 -867 46
rect -821 -200 -818 46
rect -870 -354 -818 -200
rect -634 46 -582 358
tri -289 178 -255 202 se
rect -255 178 -114 202
tri -114 178 -80 202 sw
tri -346 138 -289 178 se
rect -289 150 -80 178
rect -289 138 -255 150
tri -255 138 -238 150 nw
tri -131 138 -114 150 ne
rect -114 138 -80 150
rect -634 -200 -631 46
rect -585 -200 -582 46
rect -634 -252 -582 -200
tri -380 115 -346 138 se
rect -346 115 -289 138
tri -289 115 -255 138 nw
tri -114 115 -81 138 ne
rect -81 115 -80 138
rect -380 114 -289 115
tri -81 114 -80 115 ne
tri -80 114 10 178 sw
rect -380 88 -327 114
tri -327 88 -289 114 nw
tri -80 88 -43 114 ne
rect -43 88 10 114
rect -380 46 -328 88
rect -380 -200 -378 46
rect -332 -200 -328 46
rect -380 -252 -328 -200
rect -211 46 -159 88
rect -211 -200 -208 46
rect -162 -200 -159 46
rect -1091 -359 -963 -354
rect -1091 -405 -1045 -359
rect -999 -405 -963 -359
rect -1091 -414 -963 -405
rect -900 -355 -818 -354
rect -900 -358 -790 -355
rect -900 -410 -871 -358
rect -819 -410 -790 -358
rect -900 -414 -790 -410
rect -1434 -509 -1332 -504
rect -1434 -555 -1405 -509
rect -1359 -555 -1332 -509
rect -1434 -564 -1332 -555
rect -1211 -508 -1125 -504
rect -1211 -560 -1194 -508
rect -1142 -560 -1125 -508
rect -1211 -564 -1125 -560
rect -1070 -508 -960 -504
rect -1070 -560 -1027 -508
rect -975 -560 -960 -508
rect -1070 -564 -960 -560
rect -1027 -567 -960 -564
rect -1534 -718 -1531 -672
rect -1485 -718 -1482 -672
rect -1534 -782 -1482 -718
rect -1367 -674 -1315 -612
rect -1367 -720 -1364 -674
rect -1318 -720 -1315 -674
rect -1367 -1052 -1315 -720
rect -1027 -679 -975 -567
rect -1027 -725 -1023 -679
rect -977 -725 -975 -679
rect -1027 -782 -975 -725
rect -870 -677 -818 -414
tri -245 -490 -211 -463 se
rect -211 -488 -159 -200
rect -42 46 10 88
rect -42 -200 -38 46
rect 8 -200 10 46
rect 202 46 254 358
rect 202 -200 205 46
rect 251 -200 254 46
tri -42 -210 -41 -200 ne
rect -41 -252 10 -200
tri 10 -252 11 -200 sw
rect 202 -252 254 -200
rect 444 46 504 88
rect 444 -200 451 46
rect 497 -200 504 46
rect 444 -324 504 -200
rect 604 46 656 358
rect 604 -200 608 46
rect 654 -200 656 46
rect 604 -252 656 -200
rect 773 46 825 114
rect 773 -200 776 46
rect 822 -200 825 46
rect 444 -376 448 -324
rect 500 -376 504 -324
rect -211 -490 -162 -488
tri -162 -490 -159 -488 nw
tri 2 -490 43 -449 se
rect 43 -463 245 -449
tri 245 -463 258 -449 sw
rect 43 -490 258 -463
tri -256 -499 -245 -490 se
rect -245 -499 -173 -490
tri -173 -499 -162 -490 nw
tri -7 -499 2 -490 se
rect 2 -499 258 -490
tri 258 -499 294 -463 sw
tri -294 -530 -256 -499 se
rect -256 -530 -211 -499
tri -211 -530 -173 -499 nw
tri -30 -523 -7 -499 se
rect -7 -501 294 -499
rect -7 -523 43 -501
tri 43 -523 65 -501 nw
tri 223 -523 245 -501 ne
rect 245 -523 294 -501
tri -37 -530 -30 -523 se
rect -30 -530 21 -523
tri -313 -545 -294 -530 se
rect -294 -545 -230 -530
tri -230 -545 -211 -530 nw
tri -41 -533 -37 -530 se
rect -37 -533 21 -530
rect -41 -545 21 -533
tri 21 -545 43 -523 nw
tri 245 -536 258 -523 ne
rect 258 -536 294 -523
tri 294 -536 332 -499 sw
tri 258 -545 267 -536 ne
rect 267 -545 332 -536
tri -319 -550 -313 -545 se
rect -313 -550 -236 -545
tri -236 -550 -230 -545 nw
tri -377 -596 -319 -550 se
rect -319 -596 -294 -550
tri -294 -596 -236 -550 nw
tri -381 -600 -377 -596 se
rect -377 -600 -298 -596
tri -298 -600 -294 -596 nw
rect -870 -723 -867 -677
rect -821 -723 -818 -677
rect -870 -782 -818 -723
rect -702 -677 -650 -612
rect -702 -723 -699 -677
rect -653 -723 -650 -677
rect -702 -1052 -650 -723
rect -550 -677 -498 -612
rect -550 -723 -547 -677
rect -501 -723 -498 -677
rect -550 -857 -498 -723
rect -381 -680 -329 -600
tri -329 -625 -298 -600 nw
rect -381 -726 -378 -680
rect -332 -726 -329 -680
rect -381 -782 -329 -726
rect -41 -677 11 -545
tri 11 -555 21 -545 nw
tri 267 -555 277 -545 ne
rect 277 -555 332 -545
tri 277 -558 280 -555 ne
rect -41 -723 -38 -677
rect 8 -723 11 -677
rect -41 -780 11 -723
rect 128 -677 180 -612
rect 128 -723 131 -677
rect 177 -723 180 -677
tri 125 -835 128 -833 se
rect 128 -835 180 -723
tri -498 -857 -476 -835 sw
tri 104 -855 125 -835 se
rect 125 -855 180 -835
tri 102 -857 104 -855 se
rect 104 -857 178 -855
tri 178 -857 180 -855 nw
rect 280 -677 332 -555
rect 280 -723 283 -677
rect 329 -723 332 -677
tri -550 -931 -476 -857 ne
tri -476 -892 -441 -857 sw
tri 85 -873 102 -857 se
rect 102 -873 161 -857
tri 161 -873 178 -857 nw
tri 65 -892 85 -873 se
rect 85 -892 100 -873
rect -476 -931 100 -892
tri 100 -931 161 -873 nw
tri -476 -944 -463 -931 ne
rect -463 -944 85 -931
tri 85 -944 100 -931 nw
rect 280 -1052 332 -723
rect 444 -678 504 -376
rect 557 -329 724 -320
rect 557 -375 651 -329
rect 697 -375 724 -329
rect 557 -380 724 -375
rect 773 -490 825 -200
rect 943 46 995 358
rect 943 -200 946 46
rect 992 -200 995 46
rect 943 -252 995 -200
rect 1112 46 1164 88
rect 1112 -200 1115 46
rect 1161 -200 1164 46
rect 574 -495 684 -490
rect 574 -547 604 -495
rect 656 -547 684 -495
rect 574 -550 684 -547
rect 744 -495 854 -490
rect 744 -547 772 -495
rect 824 -547 854 -495
rect 744 -550 854 -547
rect 934 -499 1064 -490
rect 934 -545 991 -499
rect 1037 -545 1064 -499
rect 934 -550 1064 -545
rect 444 -724 451 -678
rect 497 -724 504 -678
rect 444 -782 504 -724
rect 604 -674 656 -550
rect 604 -720 608 -674
rect 654 -720 656 -674
rect 604 -782 656 -720
rect 943 -673 995 -612
rect 943 -719 946 -673
rect 992 -719 995 -673
rect 943 -1052 995 -719
rect 1112 -677 1164 -200
rect 1112 -723 1115 -677
rect 1161 -723 1164 -677
rect 1112 -782 1164 -723
rect -1599 -1074 1250 -1052
rect -1599 -1120 -1518 -1074
rect -1472 -1120 -1278 -1074
rect -1232 -1120 -1038 -1074
rect -992 -1120 -798 -1074
rect -752 -1120 -558 -1074
rect -512 -1120 -318 -1074
rect -272 -1120 -78 -1074
rect -32 -1120 162 -1074
rect 208 -1120 402 -1074
rect 448 -1120 642 -1074
rect 688 -1120 882 -1074
rect 928 -1120 1122 -1074
rect 1168 -1120 1250 -1074
rect -1599 -1192 1250 -1120
<< via1 >>
rect -871 -410 -819 -358
rect -1194 -560 -1142 -508
rect -1027 -560 -975 -508
rect 448 -376 500 -324
rect 604 -547 656 -495
rect 772 -547 824 -495
<< metal2 >>
rect 432 -319 520 -299
rect 624 -319 716 -302
rect 432 -324 716 -319
rect -1062 -354 -972 -333
rect -884 -354 -802 -341
rect -1062 -358 -802 -354
rect -1062 -410 -871 -358
rect -819 -410 -802 -358
rect 432 -376 448 -324
rect 500 -376 716 -324
rect 432 -379 716 -376
rect 432 -399 520 -379
rect 624 -402 716 -379
rect -1062 -414 -802 -410
rect -1062 -432 -972 -414
rect -884 -428 -802 -414
rect -1454 -504 -1332 -482
rect 590 -490 666 -480
rect 760 -490 835 -470
rect 964 -490 1056 -472
rect 574 -495 1056 -490
rect -1207 -504 -1127 -495
rect -1037 -504 -960 -495
rect -1454 -508 -960 -504
rect -1454 -560 -1194 -508
rect -1142 -560 -1027 -508
rect -975 -560 -960 -508
rect 574 -547 604 -495
rect 656 -547 772 -495
rect 824 -547 1056 -495
rect 574 -550 1056 -547
rect 590 -554 666 -550
rect -1454 -564 -960 -560
rect -1454 -582 -1332 -564
rect -1207 -573 -1127 -564
rect -1037 -572 -960 -564
rect 760 -566 835 -550
rect 964 -572 1056 -550
<< labels >>
rlabel nwell -1662 -417 1299 530 1 VDD
port 1 n
rlabel psubdiffcont -798 -1120 -752 -1074 1 VSS
port 2 n
rlabel polysilicon -300 -1032 914 -982 1 A
port 3 n
rlabel polysilicon -1284 288 100 338 1 B
port 4 n
rlabel metal1 -1534 -672 -1482 -200 1 L
port 5 n
rlabel metal1 -245 -530 -211 -490 1 E
port 6 n
rlabel metal1 1112 -677 1164 -200 1 G
port 7 n
<< properties >>
string path -8.850 -5.650 -8.850 2.530 -6.165 4.400 -3.060 4.400 -0.410 2.525 -0.375 -5.650 
<< end >>
