* Extracted by KLayout with GF180MCU LVS runset on : 03/10/2025 15:40

.SUBCKT gf180mcu_gp9t3v3__comp2_2 VSS A L E G B VDD
M$1 L \$22 VDD VDD pfet_03v3 L=0.3U W=3.4U AS=1.377P AD=0.918P PS=6.72U PD=4.48U
M$3 \$21 A VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U PD=4.48U
M$4 VDD B \$39 VDD pfet_03v3 L=0.3U W=3.4U AS=1.377P AD=0.918P PS=6.72U PD=4.48U
M$6 E \$27 \$39 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U
+ PD=4.48U
M$7 VDD B \$27 VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U PD=2.24U
M$8 G \$24 VDD VDD pfet_03v3 L=0.3U W=3.4U AS=0.918P AD=1.377P PS=4.48U PD=6.72U
M$10 \$22 B VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U
+ PD=2.24U
M$11 VDD \$21 \$22 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.459P PS=2.24U
+ PD=2.24U
M$12 \$39 \$21 VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.459P PS=2.24U
+ PD=2.24U
M$13 E A \$39 VDD pfet_03v3 L=0.3U W=3.4U AS=0.918P AD=1.377P PS=4.48U PD=6.72U
M$15 \$24 \$27 VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U
+ PD=2.24U
M$16 VDD A \$24 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U
+ PD=4.48U
M$17 VSS B \$27 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$18 G \$24 VSS VSS nfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.6885P PS=2.78U
+ PD=4.17U
M$20 L \$22 VSS VSS nfet_03v3 L=0.3U W=1.7U AS=0.6885P AD=0.459P PS=4.17U
+ PD=2.78U
M$22 \$21 A VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.2295P AD=0.459P PS=1.39U
+ PD=2.78U
M$23 \$35 \$27 \$24 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.102P PS=2.78U
+ PD=1.09U
M$24 VSS A \$35 VSS nfet_03v3 L=0.3U W=0.85U AS=0.102P AD=0.459P PS=1.09U
+ PD=2.78U
M$25 \$31 B VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.102P PS=2.78U
+ PD=1.09U
M$26 \$22 \$21 \$31 VSS nfet_03v3 L=0.3U W=0.85U AS=0.102P AD=0.459P PS=1.09U
+ PD=2.78U
M$27 VSS B \$23 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$28 \$26 \$27 VSS VSS nfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.6885P PS=2.78U
+ PD=4.17U
M$30 E \$21 \$23 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$31 \$26 A E VSS nfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.6885P PS=2.78U PD=4.17U
.ENDS gf180mcu_gp9t3v3__comp2_2
