VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO comp2_1x
  CLASS BLOCK ;
  FOREIGN comp2_1x ;
  ORIGIN 8.310 5.960 ;
  SIZE 14.805 BY 8.610 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -8.310 -2.085 6.495 2.650 ;
      LAYER Metal1 ;
        RECT -7.995 1.790 6.250 2.490 ;
        RECT -6.835 -1.260 -6.575 1.790 ;
        RECT -5.130 -1.260 -4.870 1.790 ;
        RECT -3.170 -1.260 -2.910 1.790 ;
        RECT 1.010 -1.260 1.270 1.790 ;
        RECT 3.020 -1.260 3.280 1.790 ;
        RECT 4.715 -1.260 4.975 1.790 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.215 -2.245 0.215 -2.505 -0.045 -2.505 ;
        RECT 0.215 -2.315 1.225 -2.245 ;
        POLYGON 1.225 -2.245 1.290 -2.315 1.225 -2.315 ;
        RECT 0.215 -2.505 1.290 -2.315 ;
        POLYGON 1.290 -2.315 1.480 -2.505 1.290 -2.505 ;
        POLYGON -0.045 -2.505 -0.045 -2.615 -0.150 -2.615 ;
        RECT -0.045 -2.615 0.055 -2.505 ;
        POLYGON -0.150 -2.615 -0.150 -2.650 -0.185 -2.650 ;
        RECT -0.150 -2.650 0.055 -2.615 ;
        POLYGON -0.185 -2.650 -0.185 -2.665 -0.205 -2.665 ;
        RECT -0.185 -2.665 0.055 -2.650 ;
        RECT -6.835 -5.260 -6.575 -3.060 ;
        RECT -3.510 -5.260 -3.250 -3.060 ;
        RECT -0.205 -3.900 0.055 -2.665 ;
        POLYGON 0.055 -2.505 0.325 -2.505 0.055 -2.775 ;
        POLYGON 1.115 -2.505 1.385 -2.505 1.385 -2.775 ;
        RECT 1.385 -2.680 1.480 -2.505 ;
        POLYGON 1.480 -2.505 1.660 -2.680 1.480 -2.680 ;
        RECT 1.385 -2.775 1.660 -2.680 ;
        POLYGON 1.385 -2.775 1.400 -2.775 1.400 -2.790 ;
        RECT 1.400 -5.260 1.660 -2.775 ;
        RECT 4.715 -5.260 4.975 -3.060 ;
        RECT -7.995 -5.960 6.250 -5.260 ;
    END
  END VSS
  PIN L
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT -7.670 -3.910 -7.410 0.440 ;
    END
  END L
  PIN E
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal1 ;
        POLYGON -1.055 -2.315 -1.055 -2.450 -1.225 -2.450 ;
        RECT -1.055 -2.440 -0.795 0.440 ;
        RECT -1.055 -2.450 -0.810 -2.440 ;
        POLYGON -0.810 -2.440 -0.795 -2.440 -0.810 -2.450 ;
        POLYGON -1.225 -2.450 -1.225 -2.495 -1.280 -2.495 ;
        RECT -1.225 -2.495 -0.865 -2.450 ;
        POLYGON -0.865 -2.450 -0.810 -2.450 -0.865 -2.495 ;
        POLYGON -1.280 -2.495 -1.280 -2.650 -1.470 -2.650 ;
        RECT -1.280 -2.650 -1.055 -2.495 ;
        POLYGON -1.055 -2.495 -0.865 -2.495 -1.055 -2.650 ;
        POLYGON -1.470 -2.650 -1.470 -2.725 -1.565 -2.725 ;
        RECT -1.470 -2.725 -1.150 -2.650 ;
        POLYGON -1.150 -2.650 -1.055 -2.650 -1.150 -2.725 ;
        POLYGON -1.565 -2.725 -1.565 -2.750 -1.595 -2.750 ;
        RECT -1.565 -2.750 -1.180 -2.725 ;
        POLYGON -1.180 -2.725 -1.150 -2.725 -1.180 -2.750 ;
        POLYGON -1.595 -2.750 -1.595 -2.980 -1.885 -2.980 ;
        RECT -1.595 -2.980 -1.470 -2.750 ;
        POLYGON -1.470 -2.750 -1.180 -2.750 -1.470 -2.980 ;
        POLYGON -1.885 -2.980 -1.885 -3.000 -1.905 -3.000 ;
        RECT -1.885 -3.000 -1.490 -2.980 ;
        POLYGON -1.490 -2.980 -1.470 -2.980 -1.490 -3.000 ;
        RECT -1.905 -3.910 -1.645 -3.000 ;
        POLYGON -1.645 -3.000 -1.490 -3.000 -1.645 -3.125 ;
    END
  END E
  PIN G
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.560 -3.910 5.820 0.440 ;
    END
  END G
  OBS
      LAYER Metal1 ;
        POLYGON -1.275 1.010 -1.275 0.890 -1.445 0.890 ;
        RECT -1.275 0.890 -0.570 1.010 ;
        POLYGON -0.570 1.010 -0.400 0.890 -0.570 0.890 ;
        POLYGON -1.445 0.890 -1.445 0.690 -1.730 0.690 ;
        RECT -1.445 0.750 -0.400 0.890 ;
        RECT -1.445 0.690 -1.275 0.750 ;
        POLYGON -1.275 0.750 -1.190 0.750 -1.275 0.690 ;
        POLYGON -0.655 0.750 -0.570 0.750 -0.570 0.690 ;
        RECT -0.570 0.690 -0.400 0.750 ;
        POLYGON -1.730 0.690 -1.730 0.575 -1.900 0.575 ;
        RECT -1.730 0.575 -1.445 0.690 ;
        POLYGON -1.445 0.690 -1.275 0.690 -1.445 0.575 ;
        POLYGON -0.570 0.690 -0.405 0.690 -0.405 0.575 ;
        RECT -0.405 0.575 -0.400 0.690 ;
        RECT -1.900 0.570 -1.445 0.575 ;
        POLYGON -0.405 0.575 -0.400 0.575 -0.400 0.570 ;
        POLYGON -0.400 0.890 0.050 0.570 -0.400 0.570 ;
        RECT -1.900 0.440 -1.635 0.570 ;
        POLYGON -1.635 0.570 -1.445 0.570 -1.635 0.440 ;
        POLYGON -0.400 0.570 -0.215 0.570 -0.215 0.440 ;
        RECT -0.215 0.440 0.050 0.570 ;
        RECT -5.965 -2.520 -5.705 0.435 ;
        RECT -4.350 -1.770 -4.090 0.440 ;
        RECT -1.900 -1.260 -1.640 0.440 ;
        RECT -0.210 -1.000 0.050 0.440 ;
        POLYGON -0.210 -1.000 -0.205 -1.000 -0.205 -1.050 ;
        RECT -0.205 -1.260 0.050 -1.000 ;
        POLYGON 0.050 -1.000 0.055 -1.260 0.050 -1.260 ;
        RECT -5.455 -2.070 -4.815 -1.770 ;
        RECT -4.500 -1.775 -4.090 -1.770 ;
        RECT -4.500 -2.070 -3.950 -1.775 ;
        RECT -7.170 -2.820 -6.660 -2.520 ;
        RECT -6.055 -2.820 -5.625 -2.520 ;
        RECT -5.350 -2.820 -4.800 -2.520 ;
        RECT -5.135 -2.835 -4.800 -2.820 ;
        RECT -5.135 -3.910 -4.875 -2.835 ;
        RECT -4.350 -3.910 -4.090 -2.070 ;
        RECT -2.750 -4.285 -2.490 -3.060 ;
        POLYGON 0.640 -4.165 0.640 -4.175 0.625 -4.175 ;
        RECT 0.640 -4.175 0.900 -3.060 ;
        RECT 2.220 -3.910 2.520 0.440 ;
        RECT 2.785 -1.900 3.620 -1.600 ;
        RECT 3.865 -2.450 4.125 0.570 ;
        RECT 2.870 -2.750 3.420 -2.450 ;
        RECT 3.720 -2.750 4.270 -2.450 ;
        RECT 4.670 -2.750 5.320 -2.450 ;
        RECT 3.020 -3.910 3.280 -2.750 ;
        POLYGON -2.490 -4.175 -2.380 -4.285 -2.490 -4.285 ;
        POLYGON 0.625 -4.175 0.625 -4.275 0.520 -4.275 ;
        RECT 0.625 -4.275 0.900 -4.175 ;
        POLYGON 0.520 -4.275 0.520 -4.285 0.510 -4.285 ;
        RECT 0.520 -4.285 0.890 -4.275 ;
        POLYGON 0.890 -4.275 0.900 -4.275 0.890 -4.285 ;
        POLYGON -2.750 -4.285 -2.380 -4.285 -2.380 -4.655 ;
        POLYGON -2.380 -4.285 -2.205 -4.460 -2.380 -4.460 ;
        POLYGON 0.510 -4.285 0.510 -4.365 0.425 -4.365 ;
        RECT 0.510 -4.365 0.805 -4.285 ;
        POLYGON 0.805 -4.285 0.890 -4.285 0.805 -4.365 ;
        POLYGON 0.425 -4.365 0.425 -4.460 0.325 -4.460 ;
        RECT 0.425 -4.460 0.500 -4.365 ;
        RECT -2.380 -4.655 0.500 -4.460 ;
        POLYGON 0.500 -4.365 0.805 -4.365 0.500 -4.655 ;
        POLYGON -2.380 -4.655 -2.315 -4.655 -2.315 -4.720 ;
        RECT -2.315 -4.720 0.425 -4.655 ;
        POLYGON 0.425 -4.655 0.500 -4.655 0.425 -4.720 ;
      LAYER Metal2 ;
        RECT 2.160 -1.595 2.600 -1.495 ;
        RECT 3.120 -1.595 3.580 -1.510 ;
        RECT -5.310 -1.770 -4.860 -1.665 ;
        RECT -4.420 -1.770 -4.010 -1.705 ;
        RECT -5.310 -2.070 -4.010 -1.770 ;
        RECT 2.160 -1.895 3.580 -1.595 ;
        RECT 2.160 -1.995 2.600 -1.895 ;
        RECT 3.120 -2.010 3.580 -1.895 ;
        RECT -5.310 -2.160 -4.860 -2.070 ;
        RECT -4.420 -2.140 -4.010 -2.070 ;
        RECT -7.270 -2.520 -6.660 -2.410 ;
        RECT 2.950 -2.450 3.330 -2.400 ;
        RECT 3.800 -2.450 4.175 -2.350 ;
        RECT 4.820 -2.450 5.280 -2.360 ;
        RECT -6.035 -2.520 -5.635 -2.475 ;
        RECT -5.185 -2.520 -4.800 -2.475 ;
        RECT -7.270 -2.820 -4.800 -2.520 ;
        RECT 2.870 -2.750 5.280 -2.450 ;
        RECT 2.950 -2.770 3.330 -2.750 ;
        RECT -7.270 -2.910 -6.660 -2.820 ;
        RECT -6.035 -2.865 -5.635 -2.820 ;
        RECT -5.185 -2.860 -4.800 -2.820 ;
        RECT 3.800 -2.830 4.175 -2.750 ;
        RECT 4.820 -2.860 5.280 -2.750 ;
  END
END comp2_1x
END LIBRARY

