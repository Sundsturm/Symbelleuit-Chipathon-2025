VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_gp9t3v3__comp2_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_gp9t3v3__comp2_1 ;
  ORIGIN 64.035 -64.415 ;
  SIZE 14.880 BY 6.350 ;
  PIN L
    ANTENNADIFFAREA 1.377000 ;
    PORT
      LAYER Metal1 ;
        RECT -63.450 67.915 -63.190 69.355 ;
        RECT -63.715 67.655 -63.190 67.915 ;
        RECT -63.715 67.310 -63.455 67.655 ;
        RECT -63.960 66.545 -63.455 67.310 ;
        RECT -63.715 66.285 -63.305 66.545 ;
        RECT -63.565 65.670 -63.305 66.285 ;
      LAYER Metal2 ;
        RECT -63.960 66.545 -63.465 67.310 ;
    END
  END L
  PIN E
    ANTENNADIFFAREA 2.295000 ;
    PORT
      LAYER Metal1 ;
        RECT -57.705 67.800 -57.165 69.355 ;
        RECT -55.185 67.800 -54.645 69.355 ;
        RECT -58.125 65.855 -57.585 66.425 ;
      LAYER Metal2 ;
        RECT -58.005 68.650 -57.165 69.355 ;
        RECT -55.185 68.650 -54.645 69.355 ;
        RECT -58.005 68.350 -54.645 68.650 ;
        RECT -58.005 67.800 -57.165 68.350 ;
        RECT -55.185 67.800 -54.645 68.350 ;
        RECT -58.005 66.425 -57.705 67.800 ;
        RECT -58.125 65.855 -57.585 66.425 ;
        RECT -58.005 65.760 -57.705 65.855 ;
    END
  END E
  PIN G
    ANTENNADIFFAREA 1.377000 ;
    PORT
      LAYER Metal1 ;
        RECT -50.005 67.915 -49.745 69.355 ;
        RECT -50.005 67.655 -49.485 67.915 ;
        RECT -49.745 67.310 -49.485 67.655 ;
        RECT -49.745 66.545 -49.230 67.310 ;
        RECT -49.885 66.285 -49.485 66.545 ;
        RECT -49.885 65.700 -49.625 66.285 ;
      LAYER Metal2 ;
        RECT -49.725 66.545 -49.230 67.310 ;
    END
  END G
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -64.035 67.205 -49.155 70.765 ;
      LAYER Metal1 ;
        RECT -63.120 69.935 -50.070 70.635 ;
        RECT -62.605 67.655 -62.345 69.935 ;
        RECT -60.925 67.655 -60.665 69.935 ;
        RECT -59.245 67.655 -58.985 69.935 ;
        RECT -56.725 67.800 -56.465 69.935 ;
        RECT -54.205 67.655 -53.945 69.935 ;
        RECT -52.525 67.655 -52.265 69.935 ;
        RECT -50.845 67.655 -50.585 69.935 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -62.725 65.115 -62.465 66.545 ;
        RECT -61.045 65.115 -60.785 66.545 ;
        RECT -55.470 65.115 -55.210 66.545 ;
        RECT -52.405 65.115 -52.145 66.545 ;
        RECT -50.725 65.115 -50.465 66.545 ;
        RECT -63.120 64.415 -50.070 65.115 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -61.770 67.565 -61.510 69.370 ;
        RECT -63.165 66.895 -62.745 67.375 ;
        RECT -61.890 66.685 -61.510 67.565 ;
        RECT -61.890 65.695 -61.630 66.685 ;
        RECT -60.085 66.545 -59.825 69.355 ;
        RECT -58.405 67.560 -58.145 69.390 ;
        RECT -55.885 67.560 -55.625 69.355 ;
        RECT -59.510 66.885 -58.725 67.310 ;
        RECT -58.405 67.300 -55.625 67.560 ;
        RECT -57.145 66.785 -54.365 67.045 ;
        RECT -54.110 66.885 -53.615 67.315 ;
        RECT -60.105 65.695 -59.265 66.545 ;
        RECT -58.830 65.615 -58.570 66.545 ;
        RECT -57.145 65.855 -56.885 66.785 ;
        RECT -56.305 65.615 -56.045 66.545 ;
        RECT -54.625 65.695 -54.365 66.785 ;
        RECT -53.365 66.545 -53.105 69.355 ;
        RECT -51.685 67.565 -51.425 69.370 ;
        RECT -51.685 66.885 -51.305 67.565 ;
        RECT -50.445 66.895 -50.025 67.400 ;
        RECT -53.925 65.695 -53.085 66.545 ;
        RECT -51.565 65.695 -51.305 66.885 ;
        RECT -58.830 65.355 -56.045 65.615 ;
      LAYER Metal2 ;
        RECT -63.165 67.375 -62.865 67.515 ;
        RECT -63.165 66.895 -62.745 67.375 ;
        RECT -61.890 67.250 -61.510 67.565 ;
        RECT -59.685 67.250 -58.545 67.310 ;
        RECT -61.890 66.950 -58.545 67.250 ;
        RECT -63.165 65.995 -62.865 66.895 ;
        RECT -61.890 66.685 -61.510 66.950 ;
        RECT -59.685 66.885 -58.545 66.950 ;
        RECT -54.110 67.185 -53.615 67.315 ;
        RECT -51.685 67.185 -51.305 67.565 ;
        RECT -50.325 67.400 -50.025 67.515 ;
        RECT -54.110 66.885 -51.305 67.185 ;
        RECT -50.445 66.895 -50.025 67.400 ;
        RECT -60.105 65.995 -59.265 66.545 ;
        RECT -63.165 65.695 -59.265 65.995 ;
        RECT -53.925 65.995 -53.085 66.545 ;
        RECT -50.325 65.995 -50.025 66.895 ;
        RECT -53.925 65.695 -50.025 65.995 ;
  END
END gf180mcu_gp9t3v3__comp2_1
END LIBRARY

