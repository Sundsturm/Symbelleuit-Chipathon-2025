** sch_path: /foss/designs/chipathon_2025/Symbelleuit-Chipathon-2025/cells/comp2/schematic/gf180mcu_gp9t3v3__comp2_2.sch
.subckt gf180mcu_gp9t3v3__comp2_2 VDD L A E G B VSS
*.PININFO L:O G:O E:O A:I B:I VDD:I VSS:I
M17 net1 NOT_A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M18 E NOT_B net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M19 net1 B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=2 m=1
M20 E A net1 VDD pfet_03v3 L=0.3u W=1.7u nf=2 m=1
M21 E NOT_A net2 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M22 net2 B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M23 E A net3 VSS nfet_03v3 L=0.3u W=0.85u nf=2 m=1
M24 net3 NOT_B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=2 m=1
M1 NOT_B B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M2 NOT_B B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M3 NOT_A A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M4 NOT_A A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M5 net5 NOT_A net4 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M6 net4 B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M7 net5 B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M8 net5 NOT_A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M9 L net5 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=2 m=1
M10 L net5 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=2 m=1
M11 net7 NOT_B net6 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M12 net6 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M13 net7 NOT_B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M14 net7 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M15 G net7 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=2 m=1
M16 G net7 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=2 m=1
.ends
