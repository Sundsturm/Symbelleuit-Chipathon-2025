magic
tech gf180mcuC
timestamp 1755577624
<< nwell >>
rect -8 63 69 127
<< nmos >>
rect 2 21 8 38
rect 19 21 25 38
rect 36 21 42 38
rect 53 21 59 38
<< pmos >>
rect 22 72 28 106
rect 33 72 39 106
<< ndiff >>
rect -8 36 2 38
rect -8 23 -6 36
rect -1 23 2 36
rect -8 21 2 23
rect 8 36 19 38
rect 8 23 11 36
rect 16 23 19 36
rect 8 21 19 23
rect 25 36 36 38
rect 25 23 28 36
rect 33 23 36 36
rect 25 21 36 23
rect 42 36 53 38
rect 42 23 45 36
rect 50 23 53 36
rect 42 21 53 23
rect 59 36 69 38
rect 59 23 62 36
rect 67 23 69 36
rect 59 21 69 23
<< pdiff >>
rect 12 104 22 106
rect 12 74 14 104
rect 19 74 22 104
rect 12 72 22 74
rect 28 72 33 106
rect 39 104 49 106
rect 39 81 42 104
rect 47 81 49 104
rect 39 72 49 81
<< ndiffc >>
rect -6 23 -1 36
rect 11 23 16 36
rect 28 23 33 36
rect 45 23 50 36
rect 62 23 67 36
<< pdiffc >>
rect 14 74 19 104
rect 42 81 47 104
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
<< polysilicon >>
rect 22 106 28 111
rect 33 106 39 111
rect 22 68 28 72
rect 19 63 28 68
rect 33 69 39 72
rect 33 67 42 69
rect 33 65 50 67
rect 33 63 42 65
rect 19 54 25 63
rect 11 52 25 54
rect 11 50 14 52
rect 2 46 14 50
rect 20 46 25 52
rect 2 44 25 46
rect 2 38 8 44
rect 19 38 25 44
rect 36 59 42 63
rect 48 62 50 65
rect 48 59 59 62
rect 36 57 59 59
rect 36 38 42 57
rect 53 38 59 57
rect 2 16 8 21
rect 19 16 25 21
rect 36 16 42 21
rect 53 16 59 21
<< polycontact >>
rect 14 46 20 52
rect 42 59 48 65
<< metal1 >>
rect -8 120 69 127
rect -8 115 11 120
rect 16 115 35 120
rect 40 115 69 120
rect -8 113 69 115
rect 14 104 19 113
rect 42 104 47 106
rect 42 79 47 81
rect 28 78 47 79
rect 14 72 19 74
rect 26 72 28 78
rect 34 74 47 78
rect 34 72 36 74
rect 28 63 33 72
rect -6 58 33 63
rect 40 59 42 65
rect 48 59 50 65
rect -6 36 -1 58
rect 12 46 14 52
rect 20 46 22 52
rect 28 48 33 58
rect 28 43 67 48
rect -6 21 -1 23
rect 11 36 16 38
rect 11 14 16 23
rect 28 36 33 43
rect 28 21 33 23
rect 45 36 50 38
rect 45 14 50 23
rect 62 36 67 43
rect 62 21 67 23
rect -8 12 69 14
rect -8 7 11 12
rect 16 7 35 12
rect 40 7 69 12
rect -8 0 69 7
<< via1 >>
rect 28 72 34 78
rect 42 59 48 65
rect 14 46 20 52
<< metal2 >>
rect 26 78 36 79
rect 26 72 28 78
rect 34 72 36 78
rect 26 71 36 72
rect 40 65 50 66
rect 40 59 42 65
rect 48 59 50 65
rect 40 58 50 59
rect 12 52 22 53
rect 12 46 14 52
rect 20 46 22 52
rect 12 45 22 46
<< labels >>
rlabel metal2 17 49 17 49 1 A
port 1 n
rlabel metal2 45 62 45 62 1 B
port 2 n
rlabel via1 31 75 31 75 1 Y
port 3 n
rlabel nsubdiffcont 13 117 13 117 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
<< end >>
