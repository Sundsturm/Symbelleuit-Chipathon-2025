  X � 	   ) � 	   )  LIB  ?z�G�{:y��0�: � 	   ) � 	   )  gf180mccu_gp9t3v3__comp2_1        ,���������   X  x   X  x���������          ,����  V����  ����d  ����d  V����  V          ,����  V����  ����T  ����T  V����  V          ,����  V����  ����D  ����D  V����  V          ,����  V����  ����4  ����4  V����  V          ,����  V����  ����$  ����$  V����  V          ,   n  V   n  �    �    V   n  V          ,  ^  V  ^  �  �  �  �  V  ^  V          ,  N  V  N  �  �  �  �  V  N  V          ,  >  V  >  �  �  �  �  V  >  V          ,���~  V���~  �     �     V���~  V          ,���^������^   X����   X����������^���          ,  ����  �   X  0   X  0���  ����          ,������������������d������d������������          ,������������������T������T������������          ,������������������D������D������������          ,������������������4������4������������          ,������������������$������$������������          ,���~�������~���   ���   �������~����          ,   n����   n���  ���  ����   n����          ,  ^����  ^���  ����  �����  ^����          ,  N����  N���  ����  �����  N����          ,  >����  >���  ����  �����  >����          ,  E���  E����  j����  j���  E���          ,   ����   �����  	����  	���   ����          ,�������������������������������������          ,���������������   �����   �����������          ,���$������$�������S�������S������$���          4   	����   	����   E����   E����   ����   	����          ,���2�������2   ����n   ����n�������2����          ,  �����  ����n  ����n  �����  �����          ,  �����  �����  �����  �����  �����          ,���������������>������>���������������          ,  �����  ����H  ����H  �����  �����          ,  Y����  Y����  �����  �����  Y����          ,������^����������n�������n���^������^          ,�������S�����������������������S�������S          ,���*���I���*���{�������{�������I���*���I          ,������������   �����   �����������������          ,���8�������8�����������������������8����          ,  ����  ����  V����  V����  ����          ,�������T���������������������T�������T          ,���a�������a���I�������I�����������a����          ,���������������I���/���I���/������������          ,���K�������K���I�������I�����������K����          ,���������������S���7���S���7������������          ,���8�������8�������t�������t�������8����          ,  ����H  �   �  �   �  ����H  ����H          ,���������������T�������T����������������          ,   �����   ����%  ����%  �����   �����          ,�������>����   ����   �������>�������>          ,  ����n  �����  \����  \���n  ����n          ,������������   �����   �����������������          ,   (���%   (   �   d   �   d���%   (���%          ,   ����      �  \   �  \����   ����          ,  �����  �   �     �  ����  �����          ,���*���{���*   ����f   ����f���{���*���{          ,�������{����   ����   �������{�������{          ,���~���{���~   �����   ��������{���~���{          ,   ����%   �   �     �  ���%   ����%          ,����   �����  ����  ����   �����   �          ,����   �����   �����   �����   �����   �          ,����   �����   �����   �����   �����   �          ,����  ����  9   d  9   d  ����            ,   (   �   (     d     d   �   (   �          ,���2   ����2   ����f   ����f   ����2   �          ,   (   �   (   �   d   �   d   �   (   �          ,���2   ����2   ����n   ����n   ����2   �          ,���*   ����*   ����f   ����f   ����*   �          ,   (   �   (   �     �     �   (   �          ,�������I�������{���/���{���/���I�������I          ,���a���I���a���{�������{�������I���a���I          ,   ���<   ���n  ����n  ����<   ���<          ,  �����  �����  V����  V����  �����          ,   	����   	���%   d���%   d����   	����          ,����������������������������������������          ,  ����  ����  V����  V����  ����          ,���8�������8�������t�������t�������8����          ,�������5�������[  V���[  V���5�������5          ,�������������������/�������/������������          ,�������������������/�������/������������          ,���a�������a����  �����  ��������a����          ,���a�������a�����������������������a����          ,�������������������/�������/������������          ,���K�������K�����������������������K����          ,�������[�����������/�������/���[�������[          ,���a�������a�����������������������a����          ,  �����  �����  �����  �����  �����          ,  ����  ����  V����  V����  ����          ,  ����  ����  V����  V����  ����          ,  ���[  ����  V����  V���[  ���[          ,�������������������7�������7������������          ,����������������������������������������          ,�������������������7�������7������������      !    ,  �����  �����  '����  '����  �����      !    ,��������������0�������0��������������      !    ,���/���w���/�������[�������[���w���/���w      !    ,���  m���  ����/  ����/  m���  m      !    ,����  m����  ����  ����  m����  m      !    ,����  m����  ����  ����  m����  m      !    ,����  m����  �����  �����  m����  m      !    ,����  m����  �����  �����  m����  m      !    ,   �  m   �  �   �  �   �  m   �  m      !    ,  �  m  �  �  �  �  �  m  �  m      !    ,  �  m  �  �  �  �  �  m  �  m      !    ,  s  m  s  �  �  �  �  m  s  m      !    ,����  m����  �����  �����  m����  m      !    ,  |���9  |���e  ����e  ����9  |���9      !    ,  |����  |����  �����  �����  |����      !    ,  |     |   -  �   -  �     |         !    ,  $���9  $���e  P���e  P���9  $���9      !    ,  $����  $����  P����  P����  $����      !    ,  $     $   -  P   -  P     $         !    ,  ����9  ����e  ���e  ���9  ����9      !    ,  �����  �����  ����  ����  �����      !    ,  �     �   -     -       �         !    ,���~   ���~   -����   -����   ���~         !    ,���~�������~�����������������������~����      !    ,���~���9���~���e�������e�������9���~���9      !    ,���>   ���>   -���j   -���j   ���>         !    ,���>�������>�������j�������j�������>����      !    ,���>���9���>���e���j���e���j���9���>���9      !    ,����   ����   -���   -���   ����         !    ,��������������������������������������      !    ,�������9�������e������e������9�������9      !    ,����   ����   -����   -����   ����         !    ,����������������������������������������      !    ,�������9�������e�������e�������9�������9      !    ,���6   ���6   -���b   -���b   ���6         !    ,���6�������6�������b�������b�������6����      !    ,���6���9���6���e���b���e���b���9���6���9      !    ,����   ����   -���
   -���
   ����         !    ,�������������������
�������
������������      !    ,�������9�������e���
���e���
���9�������9      !    ,����   ����   -����   -����   ����         !    ,����������������������������������������      !    ,�������9�������e�������e�������9�������9      !    ,���1   ���1   -���]   -���]   ���1         !    ,���1�������1�������]�������]�������1����      !    ,���1���9���1���e���]���e���]���9���1���9      !    ,����   ����   -      -      ����         !    ,����������������   ����   ������������      !    ,�������9�������e   ���e   ���9�������9      !    ,   �      �   -   �   -   �      �         !    ,   �����   �����   �����   �����   �����      !    ,   ����9   ����e   ����e   ����9   ����9      !    ,  ,     ,   -  X   -  X     ,         !    ,  ,����  ,����  X����  X����  ,����      !    ,  ,���9  ,���e  X���e  X���9  ,���9      !    ,  �     �   -     -       �         !    ,  �����  �����  ����  ����  �����      !    ,  ����9  ����e  ���e  ���9  ����9      !    ,  a���V  a����  �����  ����V  a���V      !    ,  ����R  ����~  ����~  ����R  ����R      !    ,  ���S  ���  9���  9���S  ���S      !    ,   e���S   e���   ����   ����S   e���S      !    ,�������S���������������������S�������S      !    ,�������P�������|�������|�������P�������P      !    ,�������S����������+������+���S�������S      !    ,���W���S���W�����������������S���W���S      !    ,�������S���������������������S�������S      !    ,�������V���������������������V�������V      !    ,���D���X���D�������p�������p���X���D���X      !    ,  ���S  ���  I���  I���S  ���S      !    ,  v���W  v����  �����  ����W  v���W      !    ,������Q������}���3���}���3���Q������Q      !    ,����������������/������/�����������      !    ,������������������������������������      !    ,������������������������������������      !    ,��������������������������������������      !    ,��������������������������������������      !    ,��������������������������������������      !    ,   �����   ����   ����   �����   �����      !    ,  �����  ����  ����  �����  �����      !    ,  �����  ����  ����  �����  �����      !    ,  s����  s���  ����  �����  s����      !    ,  ����  ����.  ����.  ����  ����      "    L�������������������������������F������F�������7�������7���������   	   "    !     �   �  j����  j   	   "    !     �   �����������   	   "    !     4 �������������	   	   "    !     4   �����  ����	   	   "    !     4 ���m�������m���	   	   "    !     4 4   {����   {����   R�������6������������������   	   "    !     4 $������������������L���9���L   >   	   "    !     4 �����������  M   	   "    !     4 $���r�������r���������������   >   	   "    !     4 ���T������T  _   	   "    !     4 $���[������[���:�����������   >   	   "    !     4 $������������������G���%���G   >   	   "    !     4 4���������������   ���*   ����*  #����  #����   	   "    !     4 $  3���  3���E  ����  �   >   	   "    !     4   :���  :  [   	   "    !     4   v���  v���   	   "    !     4 $   ����   �  I   �  I   �  b   	   "    !     4 $  ����  �����  B���]  B   >   	   "    !     4   ����  �  L   	   "    !     4   �   >  ����   	   "    !     4 4�����������   e���	   �����   �����   e�������   	   "    !     4 �����������  U      "    ,���E�������E���������������������E����      "    ,������^����������n�������n���^������^      "    ,������n����������������������n������n      "    ,  ���q  ����  }����  }���q  ���q      "    ,  ����n  �����  B����  B���n  ����n      "    ,���������������>������>���������������      "    ,  �����  ����H  ����H  �����  �����      "    ,  >����  >���2  ����2  �����  >����      #    ,������� �������4�������4������� �������       #    ,����������������7������7�����������      #    ,  (����  (����  \����  \����  (����      #    ,���2���r���2�������f�������f���r���2���r      #    ,���V�������V���������������������V����      #    ,���*���s���*�������^�������^���s���*���s      #    ,  �����  �����  +����  +����  �����      #    ,  \����  \���#  ����#  �����  \����      #    ,  �����  ����3  ����3  �����  �����      $    �  >����  >����  >���(  >���2  ����2  ����-  ����-  C���-  ����-  ����H  ����H  �����  �����  C����  �����  �����  �����  >����      $    l  ����n  �����  }����  }���q  ���q  ����  }����  }����  �����  �����  B����  B���n  ����n   	   $    !     < �����������(����   	   $    !     < ���7�������b����      $    ,������^����������n�������n���^������^      $    ,���������������>������>���������������          ,���^������^   X  0   X  0������^���          ,���������������2  ����2  �������������           ,����  S����  �  �  �  �  S����  S           ,���"������"����  j����  j������"���          ,�������_����  �  �  �  ����_�������_      "  
   ���W���� L       "  
     <���0 G       "  
   ���O���H E       "  
     ���� VSS       "  
       u VDD       