* SPICE3 file created from gf180mcu_gp9t3v3__comp2_1.ext - technology: gf180mcuD

X0 VDD B a_n11097_13463# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X1 a_n12405_13139# A VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X2 VSS B a_n11793_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X3 a_n10617_13139# a_n11097_13463# a_n10785_13139# VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X4 a_n10785_13139# a_n11097_13463# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X5 a_n12069_13139# B VSS VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X6 VDD a_n12633_13089# L VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X7 E a_n11097_13463# a_n11709_13531# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X8 VSS a_n12633_13089# L VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X9 a_n11457_13139# a_n11097_13463# VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X10 a_n11709_13531# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X11 E a_n12405_13139# a_n11793_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X12 G a_n10785_13139# VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X13 a_n12633_13089# a_n12405_13139# a_n12069_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X14 a_n11457_13139# A E VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X15 VSS B a_n11097_13463# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X16 E A a_n11709_13531# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X17 a_n11709_13531# a_n12405_13139# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X18 a_n12405_13139# A VDD VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X19 VDD a_n12405_13139# a_n12633_13089# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X20 VSS A a_n10617_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X21 a_n12633_13089# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X22 G a_n10785_13139# VDD VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X23 VDD A a_n10785_13139# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
C0 a_n11793_13139# a_n11457_13139# 0.20116f
C1 E a_n11457_13139# 0.12222f
C2 a_n12405_13139# VDD 0.66334f
C3 a_n11097_13463# a_n10617_13139# 0
C4 L a_n12633_13089# 0.20126f
C5 a_n12633_13089# B 0.04351f
C6 L VDD 0.21546f
C7 a_n11793_13139# a_n10785_13139# 0.00219f
C8 E a_n10785_13139# 0.01965f
C9 G B 0.00218f
C10 VDD B 1.50329f
C11 a_n11097_13463# A 0.12204f
C12 a_n10617_13139# a_n10785_13139# 0.00725f
C13 a_n12633_13089# a_n11709_13531# 0.0102f
C14 a_n11097_13463# a_n11457_13139# 0.08649f
C15 A a_n11457_13139# 0.01778f
C16 VDD a_n11709_13531# 0.44627f
C17 a_n11097_13463# a_n10785_13139# 0.48246f
C18 A a_n10785_13139# 0.04736f
C19 a_n12633_13089# a_n11793_13139# 0.09863f
C20 a_n12633_13089# E 0.03499f
C21 E G 0.00139f
C22 VDD E 0.56802f
C23 a_n11793_13139# VDD 0.00469f
C24 a_n10785_13139# a_n11457_13139# 0.11375f
C25 L a_n12405_13139# 0.01676f
C26 a_n12405_13139# B 0.11821f
C27 a_n10617_13139# VDD 0
C28 a_n11097_13463# a_n12633_13089# 0
C29 a_n12633_13089# A 0.06212f
C30 a_n11097_13463# G 0.01615f
C31 a_n12405_13139# a_n11709_13531# 0.03f
C32 a_n11097_13463# VDD 0.68777f
C33 A VDD 0.35541f
C34 a_n12633_13089# a_n11457_13139# 0.00546f
C35 VDD a_n11457_13139# 0.02145f
C36 a_n11709_13531# B 0.04739f
C37 a_n11793_13139# a_n12405_13139# 0.05556f
C38 a_n12405_13139# E 0.05439f
C39 a_n12633_13089# a_n10785_13139# 0
C40 L E 0.00125f
C41 a_n10785_13139# G 0.20881f
C42 VDD a_n10785_13139# 0.45322f
C43 E B 0.04214f
C44 a_n11793_13139# B 0.01507f
C45 a_n12633_13089# a_n12069_13139# 0.00725f
C46 a_n11097_13463# a_n12405_13139# 0.00236f
C47 A a_n12405_13139# 0.12315f
C48 a_n11793_13139# a_n11709_13531# 0.01886f
C49 E a_n11709_13531# 0.59619f
C50 a_n12069_13139# VDD 0
C51 L A 0.00223f
C52 a_n12405_13139# a_n11457_13139# 0.00828f
C53 a_n12633_13089# VDD 0.45427f
C54 a_n11097_13463# B 0.11846f
C55 A B 0.12498f
C56 VDD G 0.2164f
C57 a_n11793_13139# E 0.19862f
C58 a_n12405_13139# a_n10785_13139# 0
C59 a_n11457_13139# B 0.02796f
C60 a_n11097_13463# a_n11709_13531# 0.02399f
C61 A a_n11709_13531# 0.04833f
C62 a_n10785_13139# B 0.05942f
C63 a_n11709_13531# a_n11457_13139# 0.30402f
C64 a_n11097_13463# E 0.05504f
C65 A a_n11793_13139# 0.03927f
C66 A E 0.05261f
C67 a_n12069_13139# a_n12405_13139# 0
C68 a_n12633_13089# a_n12405_13139# 0.45949f
C69 a_n10785_13139# a_n11709_13531# 0.00623f
C70 G VSS 0.30111f
C71 E VSS 0.22261f
C72 L VSS 0.30615f
C73 VDD VSS 7.03703f
C74 a_n10617_13139# VSS 0.00558f **FLOATING
C75 a_n11457_13139# VSS 0.24f **FLOATING
C76 a_n11793_13139# VSS 0.7516f **FLOATING
C77 a_n12069_13139# VSS 0.00558f **FLOATING
C78 a_n11709_13531# VSS 0.01037f **FLOATING
C79 a_n10785_13139# VSS 0.68371f **FLOATING
C80 a_n11097_13463# VSS 0.71946f **FLOATING
C81 a_n12405_13139# VSS 0.70672f **FLOATING
C82 A VSS 1.8722f **FLOATING
C83 a_n12633_13089# VSS 0.67788f **FLOATING
C84 B VSS 0.78046f **FLOATING
