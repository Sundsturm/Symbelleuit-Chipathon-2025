  X � 	    %� 	    % LIB  >A�7KƧ�9D�/��ZT � 	    %� 	    % gf180mcu_gp9t3v3__comp2_2         ,���j ����j m��Jp m��Jp ����j �          ,��!v )��!v ���$d ���$d )��!v )          ,��!v  ����!v  �a��$d  �a��$d  ����!v  ��          ,��!v  ����!v  �a��$d  �a��$d  ����!v  ��          ,��!v )��!v ���$d ���$d )��!v )          ,��!� G��!� ���-� ���-� G��!� G          ,��8� )��8� ���;� ���;� )��8� )          ,��&& )��&& ���) ���) )��&& )          ,��=� )��=� ���@� ���@� )��=� )          ,��=� )��=� ���@� ���@� )��=� )          ,��*� )��*� ���-� ���-� )��*� )          ,��BF )��BF ���E4 ���E4 )��BF )          ,��BF )��BF ���E4 ���E4 )��BF )          ,��8� )��8� ���;� ���;� )��8� )          ,��46 )��46 ���7$ ���7$ )��46 )          ,��/� )��/� ���2t ���2t )��/� )          ,��*� )��*� ���-� ���-� )��*� )          ,��&& )��&& ���) ���) )��&& )          ,��/� )��/� ���2t ���2t )��/� )          ,��8� G��8� ���D� ���D� G��8� G          ,��.� G��.� ���7� ���7� G��.� G          ,��46 )��46 ���7$ ���7$ )��46 )          ,��BF )��BF ���E4 ���E4 )��BF )          ,��BF )��BF ���E4 ���E4 )��BF )          ,��F� )��F� ���I� ���I� )��F� )          ,��F� )��F� ���I� ���I� )��F� )          ,��F� )��F� ���I� ���I� )��F� )          ,��F� )��F� ���I� ���I� )��F� )          ,��
 )��
 ���� ���� )��
 )          ,��
 )��
 ���� ���� )��
 )          ,��� )��� ���� ���� )��� )          ,�� )�� ��� ��� )�� )          ,��f )��f ���T ���T )��f )          ,��� )��� ���� ���� )��� )          ,��
 )��
 ���� ���� )��
 )          ,�� � )�� � ���� ���� )�� � )          ,��V )��V ���D ���D )��V )          ,��� )��� ���� ���� )��� )          ,��
 )��
 ���� ���� )��
 )          ,�� G�� ��� ��� G�� G          ,��/ G��/ ��� � ��� � G��/ G          ,��� )��� ���� ���� )��� )          ,��V )��V ���D ���D )��V )          ,��f )��f ���T ���T )��f )          ,�� � )�� � ���� ���� )�� � )          ,���� )���� ����� ����� )���� )          ,���� )���� ����� ����� )���� )          ,��f  ����f  �a��T  �a��T  ����f  ��          ,���  �����  �a���  �a���  �����  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,�� �  ��� � ���� ����  ��� �  �          ,���  �����  �a���  �a���  �����  ��          ,��  ����  �a��  �a��  ����  ��          ,��f  ����f  �a��T  �a��T  ����f  ��          ,���  �����  �a���  �a���  �����  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,��V  ����V  �a��D  �a��D  ����V  ��          ,���  ���� ���7 ���7  ����  �          ,��c  ���c ���"W ���"W  ���c  �          ,��
  ����
  �a���  �a���  ����
  ��          ,���  �����  �a���  �a���  �����  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,�� �  ���� �  �a���  �a���  ���� �  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,����  ������  �a����  �a����  ������  ��          ,��/�  ����/�  �a��2t  �a��2t  ����/�  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��BF  ����BF  �a��E4  �a��E4  ����BF  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��F�  ����F�  �a��I�  �a��I�  ����F�  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��9O  ���9O ���EC ���EC  ���9O  �          ,��0�  ���0� ���8# ���8#  ���0�  �          ,��#�  ���#� ���/w ���/w  ���#�  �          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��=�  ����=�  �a��@�  �a��@�  ����=�  ��          ,��46  ����46  �a��7$  �a��7$  ����46  ��          ,��8�  ����8�  �a��;�  �a��;�  ����8�  ��          ,��8�  ����8�  �a��;�  �a��;�  ����8�  ��          ,��46  ����46  �a��7$  �a��7$  ����46  ��          ,��/�  ����/�  �a��2t  �a��2t  ����/�  ��          ,��*�  ����*�  �a��-�  �a��-�  ����*�  ��          ,��&&  ����&&  �a��)  �a��)  ����&&  ��          ,��&&  ����&&  �a��)  �a��)  ����&&  ��          ,��*�  ����*�  �a��-�  �a��-�  ����*�  ��           ,��	� ��	� �� �� ��	�            ,��� ��� ��� ��� ���            ,��R ��R ��h ��h ��R            ,��� ��� ��� ��� ���            ,�� � �� � ��� ��� �� �            ,��!b ��!b ��$x ��$x ��!b            ,��& ��& ��)( ��)( ��&            ,��*� ��*� ��-� ��-� ��*�            ,��/r ��/r ��2� ��2� ��/r            ,��4" ��4" ��78 ��78 ��4"            ,��8� ��8� ��;� ��;� ��8�            ,�� ��� ���U ���U ��� �           ,��� ���� ��� ��� ���� �           ,��� ���� ���!! ���!! ���� �           ,��  ����  ����U  ����U  ����  ��           ,���  �����  ����  ����  �����  ��           ,���  �����  ����!!  ����!!  �����  ��           ,��V ��V ��X ��X ��V            ,��=� ��=� ��@� ��@� ��=�            ,��	� ��	� �� �� ��	�            ,��	� ��	� �� �� ��	�            ,��=� ��=� ��@� ��@� ��=�            ,��V ��V ��X ��X ��V            ,���  �����  ����!!  ����!!  �����  ��           ,���  �����  ����  ����  �����  ��           ,��  ����  ����U  ����U  ����  ��           ,��� ���� ���!! ���!! ���� �           ,��� ���� ��� ��� ���� �           ,�� ��� ���U ���U ��� �           ,��8� ��8� ��;� ��;� ��8�            ,��4" ��4" ��78 ��78 ��4"            ,��/r ��/r ��2� ��2� ��/r            ,��*� ��*� ��-� ��-� ��*�            ,��& ��& ��)( ��)( ��&            ,��!b ��!b ��$x ��$x ��!b            ,��� ��� ��� ��� ���            ,�� �� �� �� ��            ,��R ��R ��h ��h ��R            ,��� ��� ��� ��� ���            ,��	� ��	� �� �� ��	�            ,���� ���� m��I� m��I� ����            ,��B2 ��B2 ��E4 ��E4 ��B2            ,��B2 ��B2 ��E4 ��E4 ��B2            ,��$� ���$� ���.A ���.A ���$� �           ,��1� ���1� ���6� ���6� ���1� �           ,��:� ���:� ���@� ���@� ���:� �           ,��$�  ����$�  ����.A  ����.A  ����$�  ��           ,��1�  ����1�  ����6�  ����6�  ����1�  ��           ,��:�  ����:�  ����@�  ����@�  ����:�  ��           ,��:�  ����:�  ����@�  ����@�  ����:�  ��           ,��1�  ����1�  ����6�  ����6�  ����1�  ��           ,��$�  ����$�  ����.A  ����.A  ����$�  ��           ,����  ������ ���E� ���E�  ������  ��           ,��:� ���:� ���@� ���@� ���:� �           ,��1� ���1� ���6� ���6� ���1� �           ,��$� ���$� ���.A ���.A ���$� �           ,��B2 ��B2 ��E4 ��E4 ��B2            ,��B2 ��B2 ��E4 ��E4 ��B2            ,��F� ��F� ��I� ��I� ��F�            ,��F� ��F� ��I� ��I� ��F�            ,��F� ��F� ��I� ��I� ��F�            ,��F� ��F� ��I� ��I� ��F�            ,�� � �� � ��� ��� �� �            ,���� ���� ���� ���� ����            ,���� ���� ���� ���� ����           ,��� ���� ���} ���} ���� �          ,��� a��� ��� ��� a��� a          ,��� a��� ���} ���} a��� a          ,���  �����  �u���  �u���  �����  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,��R  ����R  �u��h  �u��h  ����R  ��          ,��  ����  �u��  �u��  ����  ��          ,���  �����  �u���  �u���  �����  ��          ,��!b  ����!b  �u��$x  �u��$x  ����!b  ��          ,��&  ����&  �u��)(  �u��)(  ����&  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��          ,��/r  ����/r  �u��2�  �u��2�  ����/r  ��          ,��4"  ����4"  �u��78  �u��78  ����4"  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��	�  ����	�  �u��  �u��  ����	�  ��          ,��B  ����B  �u��X  �u��X  ����B  ��          ,��B  ����B  �u��X  �u��X  ����B  ��          ,��	�  ����	�  �u��  �u��  ����	�  ��          ,��8�  ����8�  �u��;�  �u��;�  ����8�  ��          ,��4"  ����4"  �u��78  �u��78  ����4"  ��          ,��/r  ����/r  �u��2�  �u��2�  ����/r  ��          ,��*�  ����*�  �u��-�  �u��-�  ����*�  ��          ,��&  ����&  �u��)(  �u��)(  ����&  ��          ,��!b  ����!b  �u��$x  �u��$x  ����!b  ��          ,���  �����  �u���  �u���  �����  ��          ,��  ����  �u��  �u��  ����  ��          ,��R  ����R  �u��h  �u��h  ����R  ��          ,��=�  ����=�  �u��@�  �u��@�  ����=�  ��          ,���  �����  �u���  �u���  �����  ��          ,��� a��� ���} ���} a��� a          ,��� a��� ��� ��� a��� a          ,��� ���� ���} ���} ���� �          ,��E ���E ���� ���� ���E �          ,��# ���# ���,� ���,� ���# �          ,��05 ���05 ���6u ���6u ���05 �          ,��: ���: ���@M ���@M ���: �          ,��# a��# ���,� ���,� a��# a          ,��05 a��05 ���6u ���6u a��05 a          ,��: a��: ���@M ���@M a��: a          ,��: a��: ���@M ���@M a��: a          ,��05 a��05 ���6u ���6u a��05 a          ,��# a��# ���,� ���,� a��# a          ,�� o ��� o ���Ek ���Ek ��� o �          ,��: ���: ���@M ���@M ���: �          ,��05 ���05 ���6u ���6u ���05 �          ,��# ���# ���,� ���,� ���# �          ,��BF  ����BF  �u��EH  �u��EH  ����BF  ��          ,��BF  ����BF  �u��EH  �u��EH  ����BF  ��          ,��BF  ����BF  �u��EH  �u��EH  ����BF  ��          ,��BF  ����BF  �u��EH  �u��EH  ����BF  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,��F�  ����F�  �u��I�  �u��I�  ����F�  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,�� �  ���� �  �u���  �u���  ���� �  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,����  ������  �u����  �u����  ������  ��          ,��K ���K ���< ���< ���K �          ,��s ���s ���� ���� ���s �          ,��	� ��	� ���
� ���
� ��	�           ,��>� U��>� ��C' ��C' U��>� U          ,��K ���K ���w ���w ���K �          ,��	C U��	C ��
� ��
� U��	C U          ,��� ���� ���w ���w ���� �          ,���  ����� ���� ����  �����  ��          ,��� ���� ���� ���� ���� �          ,��# ��# ���O ���O ��#           ,��O ��O ��� ; ��� ; ��O           ,���  ����� }�� }��  �����  ��          ,��� }��� E��� E��� }��� }          ,��� U��� �� �� U��� U          ,���  ����� U��� U���  �����  ��          ,��(� U��(� ��3� ��3� U��(� U          ,��%' ��%' ���(o ���(o ��%'           ,��:� E��:� ���< ���< E��:� E          ,��A�  ����A� U��C' U��C'  ����A�  ��          ,��>; ��>; ���B� ���B� ��>;           ,��	C  ����	C  ����6  ����6  ����	C  ��          ,��A� ���A� ���B� ���B� ���A� �          ,��	C  ����	C  ����6  ����6  ����	C  ��          ,��:� E��:� ���< ���< E��:� E          ,��4�  ����4� ��6 ��6  ����4�  ��          ,��%�  ����%� U��&� U��&�  ����%�  ��          ,��#� U��#� ��&� ��&� U��#� U          ,��#� ��#� ���%' ���%' ��#�           ,��  ���� �� ; �� ;  ����  ��          ,��  ���� }��� }���  ����  ��          ,���  ����� }�� }��  �����  ��          ,��� E��� ��� ��� E��� E          ,��k ���k ���� ���� ���k �          ,��� ���� ��� ��� ���� �          ,��� ���� ���� ���� ���� �          ,���  ����� ���� ����  �����  ��          ,��	C  ����	C U��
o U��
o  ����	C  ��          ,��� ���� ���w ���w ���� �          ,��K ���K ���w ���w ���K �          ,���  ����� U��' U��'  �����  ��          ,��� ��� ��� ��� ���           ,��s ���s ���� ���� ���s �          ,��K ���K ���< ���< ���K �          ,��+ ��+ ���� ���� ��+           ,��+ ���+ ���W ���W ���+ �          ,���  ����� U��� U���  �����  ��          ,��� U��� ��' ��' U��� U          ,��(�  ����(� U��* U��*  ����(�  ��          ,��>; ���>; ���?g ���?g ���>; �          ,��>; ��>; ��?� ��?� ��>;           ,��:� }��:� E��<� E��<� }��:� }          ,��;k  ����;k }��<� }��<�  ����;k  ��          ,��>�  ����>� U��?� U��?�  ����>�  ��          ,��;k  ����;k }��<� }��<�  ����;k  ��          ,��:� }��:� E��<� E��<� }��:� }          ,��2�  ����2� U��3� U��3�  ����2�  ��          ,��,/  ����,/ U��-[ U��-[  ����,/  ��          ,��/� ��/� ��1� ��1� ��/�           ,��4c ��4c ���6 ���6 ��4c           ,��4c ���4c ���5� ���5� ���4c �          ,��*� ��*� ���2G ���2G ��*�           ,��1 ���1 ���2G ���2G ���1 �          ,��*� ���*� ���+� ���+� ���*� �          ,��'C ���'C ���(o ���(o ���'C �      !    ,��" ���" x��#[ x��#[ ���" �      !    ,��"  ���"  ����#[  ����#[  ���"  �      !    ,��"  ���"  ����#[  ����#[  ���"  �      !    ,��" 	U��" 
1��#[ 
1��#[ 	U��" 	U      !    ,��" +��" ��#[ ��#[ +��" +      !    ,��" ��" ���#[ ���#[ ��"       !    ,��" ���" x��#[ x��#[ ���" �      !    ,��%� ��%� ���&� ���&� ��%�       !    ,��%� +��%� ��&� ��&� +��%� +      !    ,��%� 	U��%� 
1��&� 
1��&� 	U��%� 	U      !    ,��+� ���+� x��,� x��,� ���+� �      !    ,��) +��) ��)� ��)� +��) +      !    ,��0� ���0� x��1k x��1k ���0� �      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��5? ���5? x��6 x��6 ���5? �      !    ,��>� ���>� x��?{ x��?{ ���>� �      !    ,��) 	U��) 
1��)� 
1��)� 	U��) 	U      !    ,��0� ���0� x��1k x��1k ���0� �      !    ,��) +��) ��)� ��)� +��) +      !    ,��+� ���+� x��,� x��,� ���+� �      !    ,��) ��) ���)� ���)� ��)       !    ,��'/ ���'/ x��( x��( ���'/ �      !    ,��9� ���9� x��:� x��:� ���9� �      !    ,��9� ���9� x��:� x��:� ���9� �      !    ,��'/ ���'/ x��( x��( ���'/ �      !    ,��) ��) ���)� ���)� ��)       !    ,��>� ���>� x��?{ x��?{ ���>� �      !    ,��5? ���5? x��6 x��6 ���5? �      !    ,��CO ���CO x��D+ x��D+ ���CO �      !    ,��CO ���CO x��D+ x��D+ ���CO �      !    ,��CO ���CO x��D+ x��D+ ���CO �      !    ,��CO ���CO x��D+ x��D+ ���CO �      !    ,��G� ���G� x��H� x��H� ���G� �      !    ,��G� ���G� x��H� x��H� ���G� �      !    ,��G� ���G� x��H� x��H� ���G� �      !    ,��G� ���G� x��H� x��H� ���G� �      !    ,��CO 	U��CO 
1��D+ 
1��D+ 	U��CO 	U      !    ,��CO ��CO ���D+ ���D+ ��CO       !    ,��CO +��CO ��D+ ��D+ +��CO +      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��@ 	U��@ 
1��@� 
1��@� 	U��@ 	U      !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��2� ��2� ���3� ���3� ��2�       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��<� ��<� ���=� ���=� ��<�       !    ,��@ ��@ ���@� ���@� ��@       !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��@ +��@ ��@� ��@� +��@ +      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��@ 	U��@ 
1��@� 
1��@� 	U��@ 	U      !    ,��<� 	U��<� 
1��=� 
1��=� 	U��<� 	U      !    ,��9w 	U��9w 
1��:S 
1��:S 	U��9w 	U      !    ,��6/ 	U��6/ 
1��7 
1��7 	U��6/ 	U      !    ,��2� 	U��2� 
1��3� 
1��3� 	U��2� 	U      !    ,��/� 	U��/� 
1��0{ 
1��0{ 	U��/� 	U      !    ,��,W 	U��,W 
1��-3 
1��-3 	U��,W 	U      !    ,��@ +��@ ��@� ��@� +��@ +      !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��@ ��@ ���@� ���@� ��@       !    ,��<� ��<� ���=� ���=� ��<�       !    ,��9w ��9w ���:S ���:S ��9w       !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��2� ��2� ���3� ���3� ��2�       !    ,�� ��� x��� x��� ��� �      !    ,��7 +��7 ��  ��  +��7 +      !    ,�� �� ���� ���� ��       !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� ��� ���� ���� ���       !    ,��7 ��7 ���  ���  ��7       !    ,��� ���� x��� x��� ���� �      !    ,��o ���o x��K x��K ���o �      !    ,�� ��� x��� x��� ��� �      !    ,��� ���� x��� x��� ���� �      !    ,��� +��� ��� ��� +��� +      !    ,��� ��� ���� ���� ���       !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��� ���� x��� x��� ���� �      !    ,��� ���� x��� x��� ���� �      !    ,���� ����� x���� x���� ����� �      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��� ��� ���� ���� ���       !    ,��? ��? ���	 ���	 ��?       !    ,��� ��� ���c ���c ���       !    ,��� ��� ���� ���� ���       !    ,��� +��� ��� ��� +��� +      !    ,��? +��? ��	 ��	 +��? +      !    ,��� +��� ��c ��c +��� +      !    ,��� +��� ��� ��� +��� +      !    ,�� +�� ��� ��� +�� +      !    ,�� ��� x��� x��� ��� �      !    ,��� +��� ��� ��� +��� +      !    ,��_ ���_ x��; x��; ���_ �      !    ,�� ��� x��� x��� ��� �      !    ,�� +�� ��� ��� +�� +      !    ,��_ +��_ ��; ��; +��_ +      !    ,��� +��� ��c ��c +��� +      !    ,��? +��? ��	 ��	 +��? +      !    ,��� +��� ��� ��� +��� +      !    ,��_ ��_ ���; ���; ��_       !    ,��� ��� ���c ���c ���       !    ,��? ��? ���	 ���	 ��?       !    ,��� ��� ���� ���� ���       !    ,��7 	U��7 
1��  
1��  	U��7 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� 	U�� 
1��� 
1��� 	U�� 	U      !    ,��_ 	U��_ 
1��; 
1��; 	U��_ 	U      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,��� 	U��� 
1��� 
1��� 	U��� 	U      !    ,�� ��� x��� x��� ��� �      !    ,��� ���� x��� x��� ���� �      !    ,�� ��� x��� x��� ��� �      !    ,��o ���o x��K x��K ���o �      !    ,��� ���� x��� x��� ���� �      !    ,��7 ��7 ���  ���  ��7       !    ,��� ��� ���� ���� ���       !    ,��? 	U��? 
1��	 
1��	 	U��? 	U      !    ,�� �� ���� ���� ��       !    ,��7 +��7 ��  ��  +��7 +      !    ,��� 	U��� 
1��c 
1��c 	U��� 	U      !    ,��_ ���_ x��; x��; ���_ �      !    ,��� +��� ��� ��� +��� +      !    ,���� ����� x���� x���� ����� �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,��� ���� ���o ���o ���� �      !    ,��K ���K ���' ���' ���K �      !    ,�� � ��� � ���!� ���!� ��� � �      !    ,��� ���� ���� ���� ���� �      !    ,��W ���W ���3 ���3 ���W �      !    ,�� ��� ���� ���� ��� �      !    ,��  ���  �����  �����  ���  �      !    ,���  ����  �����  �����  ����  �      !    ,��_ ���_ ���; ���; ���_ �      !    ,��  ���  �����  �����  ���  �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,�� ��� ���[ ���[ ��� �      !    ,��� ���� ���� ���� ���� �      !    ,��  ���  �����  �����  ���  �      !    ,�� ��� ���� ���� ��� �      !    ,��W ���W ���3 ���3 ���W �      !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��7 ���7 ��� ��� ���7 �      !    ,���  ����  �����  �����  ����  �      !    ,��o  ���o  ����K  ����K  ���o  �      !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���[ ���[ ��� �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��� ���� ���o ���o ���� �      !    ,��_  ���_  ����;  ����;  ���_  �      !    ,��  ���  �����  �����  ���  �      !    ,��_ ���_ ���; ���; ���_ �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,��o  ���o  ����K  ����K  ���o  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,���  ����  �����  �����  ����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,����  �����  ������  ������  �����  �      !    ,��_ ���_ ���; ���; ���_ �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��1C ���1C ���2 ���2 ���1C �      !    ,��C� ���C� ���D� ���D� ���C� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��9� ���9� ���:� ���:� ���9� �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��@ ���@ ���A[ ���A[ ���@ �      !    ,��0v ���0v ���1R ���1R ���0v �      !    ,��>� ���>� ���?{ ���?{ ���>� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��1C ���1C ���2 ���2 ���1C �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��>� ���>� ���?{ ���?{ ���>� �      !    ,��0v ���0v ���1R ���1R ���0v �      !    ,��@ ���@ ���A[ ���A[ ���@ �      !    ,��'k ���'k ���(G ���(G ���'k �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��CO  ���CO  ����D+  ����D+  ���CO  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��G�  ���G�  ����H�  ����H�  ���G�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��'/  ���'/  ����(  ����(  ���'/  �      !    ,��+�  ���+�  ����,�  ����,�  ���+�  �      !    ,��0�  ���0�  ����1k  ����1k  ���0�  �      !    ,��5?  ���5?  ����6  ����6  ���5?  �      !    ,��9�  ���9�  ����:�  ����:�  ���9�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��>�  ���>�  ����?{  ����?{  ���>�  �      !    ,��9�  ���9�  ����:�  ����:�  ���9�  �      !    ,��5?  ���5?  ����6  ����6  ���5?  �      !    ,��0�  ���0�  ����1k  ����1k  ���0�  �      !    ,��+�  ���+�  ����,�  ����,�  ���+�  �      !    ,��'/  ���'/  ����(  ����(  ���'/  �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��9� ���9� ���:� ���:� ���9� �      "    ,��� ���� G��� G��� ���� �      "    ,�� ��� ��� ��� ��� �      "    ,��%� ���%� ���&� ���&� ���%� �      "    ,��� ���� ���)� ���)� ���� �      "    ,��� :��� V��� V��� :��� :      "    ,���j  �����j  �[��Jp  �[��Jp  �����j  ��      "    ,���  �K���  O��%  O��%  �K���  �K      "    ,��� ���� ���)� ���)� ���� �      "    ,��# ���# ��� ' ��� ' ���# �      "    ,�� ��� ��� ��� ��� �      "    ,��� /��� G��� G��� /��� /      "    ,���j ����j m��Jp m��Jp ����j �      "    ,��(� ���(� ���)� ���)� ���(� �      "    ,��(� ���(� ���)� ���)� ���(� �      "    ,��� E��� ���� ���� E��� E      "    ,��� ���� ��� ��� ���� �      "    ,��n ���n ���r ���r ���n �      "    ,��n ���n ���r ���r ���n �      "    ,��/� G��/� /��0� /��0� G��/� G      "    ,��C; G��C; ���D? ���D? G��C; G      "    ,��6 G��6 /��7 /��7 G��6 G      "    ,��6 G��6 ���7 ���7 G��6 G      "    ,��<� G��<� ���=� ���=� G��<� G      "    ,��/� G��/� ���0� ���0� G��/� G      "    ,��"k ���"k ���#o ���#o ���"k �      "    ,�� ; :�� ; V��"W V��"W :�� ; :      "    ,��� 	K��� ���� ���� 	K��� 	K      "    ,��� G��� ���� ���� G��� G      "    ,��� G��� ���� ���� G��� G      "    ,��O ���O ���k ���k ���O �      "    ,��K G��K ���O ���O G��K G      "    ,��+ G��+ ���	/ ���	/ G��+ G      "    ,��� G��� 	K��� 	K��� G��� G      "    ,��� 	K��� ���� ���� 	K��� 	K      "    ,��� G��� 	K��� 	K��� G��� G      "    ,��
� }��
� ���r ���r }��
� }      "    ,��
� }��
� ���r ���r }��
� }      "    ,���  �[��� ���� ����  �[���  �[      "    ,��
�  ���
� }��� }���  ���
�  �      "    ,��� O��� /��� /��� O��� O      "    ,��� ���� O��� O��� ���� �      "    ,���  �[��� ���� ����  �[���  �[      "    ,��
�  ���
� }��� }���  ���
�  �      "    ,��k  ���k ���o ���o  ���k  �      "    ,��� ���� ���o ���o ���� �      "    ,��k  ���k ���o ���o  ���k  �      "    ,��� O��� /��� /��� O��� O      "    ,��� O��� /��� /��� O��� O      "    ,��C  �[��C ���G ���G  �[��C  �[      "    ,�� ?�� ���� ���� ?�� ?      "    ,���  O��� ���� ����  O���  O      "    ,���  ���� ���7 ���7  ����  �      "    ,��'W  �[��'W ���([ ���([  �[��'W  �[      "    ,���  ���� ���7 ���7  ����  �      "    ,��#  �[��# ���' ���'  �[��#  �[      "    ,��6�  �[��6� ���7� ���7�  �[��6�  �[      "    ,��-�  �[��-� ���.� ���.�  �[��-�  �[      "    ,��=#  �[��=# ���>' ���>'  �[��=#  �[      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��$  O��$ ���% ���%  O��$  O      "    ,��=#  �[��=# ���>' ���>'  �[��=#  �[      "    ,��C�  �[��C� ���D� ���D�  �[��C�  �[      "    ,��/� E��/� ���1� ���1� E��/� E      "    ,��@k ���@k ���A� ���A� ���@k �      "    ,��@k  ���@k ���Ao ���Ao  ���@k  �      "    ,��/� E��/� ���1� ���1� E��/� E      "    ,��@k  ���@k ���Ao ���Ao  ���@k  �      "    ,��@k ���@k ���A� ���A� ���@k �      "    ,��@� ���@� O��A� O��A� ���@� �      "    ,��9�  ���9� E��:� E��:�  ���9�  �      "    ,��0�  ���0� ���3� ���3�  ���0�  �      "    ,��*�  ���*� ���+� ���+�  ���*�  �      "    ,��>; O��>; H��?� H��?� O��>; O      "    ,��>; O��>; H��?� H��?� O��>; O      "    ,��0�  ���0� ���3� ���3�  ���0�  �      "    ,��9�  ���9� E��:� E��:�  ���9�  �      "    ,��@� O��@� H��B� H��B� O��@� O      "    ,��9c E��9c ���:� ���:� E��9c E      "    ,��9c E��9c ���:� ���:� E��9c E      "    ,��+� ���+� ���-� ���-� ���+� �      "    ,��?� G��?� 	K��A� 	K��A� G��?� G      "    ,��?� 	K��?� ���@� ���@� 	K��?� 	K      "    ,��?� G��?� 	K��A� 	K��A� G��?� G      "    ,��?� 	K��?� ���@� ���@� 	K��?� 	K      "    ,��+� ���+� ���-� ���-� ���+� �      "    ,��9c ���9c ���:g ���:g ���9c �      "    ,��9c ���9c ���:g ���:g ���9c �      "    ,��2� ���2� ���3� ���3� ���2� �      "    ,��@� H��@� G��A� G��A� H��@� H      "    ,��2� ���2� ���3� ���3� ���2� �      "    ,�� ��� ���+� ���+� ��� �      #    ,��� ��� ��� ��� ���       #    ,��� 
��� ��� ��� 
��� 
      #    ,��X ���X ���\ ���\ ���X �      #    ,��K ���K ���O ���O ���K �      #    ,��- ��- ��1 ��1 ��-       #    ,�� � ��� � ���!� ���!� ��� � �      #    ,��: ���: ���> ���> ���: �      #    ,��K ���K ���O ���O ���K �      #    ,��7 ���7 ���; ���; ���7 �      #    ,��- ��- ��1 ��1 ��-       #    ,��K ���K ���O ���O ���K �      #    ,��X ���X ���\ ���\ ���X �      #    ,��,C ��,C ��-G ��-G ��,C       #    ,��,C 
��,C ��-G ��-G 
��,C 
      #    ,��0b ���0b ���1f ���1f ���0b �      #    ,��9� ��9� ��:� ��:� ��9�       #    ,��>� ���>� ���?� ���?� ���>� �      #    ,��A� ���A� ���B� ���B� ���A� �      #    ,��2y ���2y ���3} ���3} ���2y �      #    ,��2y ���2y ���3} ���3} ���2y �      #    ,��A� ���A� ���B� ���B� ���A� �      #    ,��>� ���>� ���?� ���?� ���>� �      #    ,��9� ��9� ��:� ��:� ��9�       #    ,��0b ���0b ���1f ���1f ���0b �      #    ,��,C 
��,C ��-G ��-G 
��,C 
      #    ,��,C ��,C ��-G ��-G ��,C       $    ,��� E��� ���� ���� E��� E      $    ,��/� E��/� q��:� q��:� E��/� E      $    ,��� O��� /��� /��� O��� O      $    ,��
� ���
� ���r ���r ���
� �      $    ,��� :��� V��� V��� :��� :      $    ,�� ; :�� ; V��"W V��"W :�� ; :      $    ,��� ���� O��' O��' ���� �      $    ,��
� }��
� ���r ���r }��
� }      $    ,��� :��� V��"W V��"W :��� :      $    ,��� ���� ���7 ���7 ���� �      $    ,���  ���� ���7 ���7  ����  �      $    ,���  ���� ���7 ���7  ����  �      $    ,��� ���� ���7 ���7 ���� �      $    ,��
� }��
� ���r ���r }��
� }      $    ,��� ���� O��' O��' ���� �      $    ,��
� ���
� ��� ��� ���
� �      $    ,��
� ���
� ���r ���r ���
� �      $    ,��� O��� /��� /��� O��� O      $    ,��� O��� /��� /��� O��� O      $    ,��� /��� ���� ���� /��� /      $    ,��O V��O 
���k 
���k V��O V      $    ,��O *��O ���k ���k *��O *      $    ,��+� *��+� ���-� ���-� *��+� *      $    ,��+� ���+� 
���-� 
���-� ���+� �      $    ,��/� q��/� ���1� ���1� q��/� q      $    ,��9c q��9c ���:� ���:� q��9c q      $    ,��>� H��>� ���?� ���?� H��>� H      $    ,��>; O��>; H��?� H��?� O��>; O      $    ,��0� ���0� ���3� ���3� ���0� �      $    ,��>� ���>� O��?� O��?� ���>� �      $    ,��0�  ���0� ���?� ���?�  ���0�  �      $    ,��0�  ���0� ���?� ���?�  ���0�  �      $    ,��@� O��@� H��B� H��B� O��@� O      $    ,��>� ���>� O��?� O��?� ���>� �      $    ,��0� ���0� ���3� ���3� ���0� �      $    ,��>; O��>; H��?� H��?� O��>; O      $    ,��/� |��/� ���:� ���:� |��/� |      $    ,��>� H��>� ���?� ���?� H��>� H      $    ,��9c q��9c ���:� ���:� q��9c q      $    ,��/� q��/� ���1� ���1� q��/� q      $    ,��+� ���+� 
���-� 
���-� ���+� �      $    ,��O 
���O *��-� *��-� 
���O 
�      $    ,��+� *��+� ���-� ���-� *��+� *      $  
      @Y������ ��AL | G       $  
      @Y������ ��� : L       $  
      @Y������ ��� J E       "  
      @I�^5?|� ��7�  VDD       "  
      @I�^5?|� ��7�  �� VSS         
 ��
V � A         
 ��� � B         
 ��� � B         
 ��
V � A       