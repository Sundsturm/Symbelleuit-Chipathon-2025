* NGSPICE file created from gf180mcu_gp9t3v3__comp2_1.ext - technology: gf180mcuD

.subckt gf180mcu_gp9t3v3__comp2_1 VDD L A E G B VSS
X0 VDD.t7 B.t0 a_n11097_13463# VDD.t6 pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X1 a_n12405_13139# A.t0 VSS.t15 VSS.t14 nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X2 VSS.t7 B.t1 a_n11793_13139# VSS.t6 nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X3 a_n10617_13139# a_n11097_13463# a_n10785_13139# VSS.t10 nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X4 a_n10785_13139# a_n11097_13463# VDD.t10 VDD.t9 pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X5 a_n12069_13139# B.t2 VSS.t5 VSS.t4 nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X6 VDD.t21 a_n12633_13089# L.t1 VDD.t20 pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X7 E.t0 a_n11097_13463# a_n11709_13531# VDD.t8 pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X8 VSS.t19 a_n12633_13089# L.t0 VSS.t18 nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X9 a_n11457_13139# a_n11097_13463# VSS.t9 VSS.t8 nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X10 a_n11709_13531# B.t3 VDD.t5 VDD.t4 pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X11 E.t3 a_n12405_13139# a_n11793_13139# VSS.t17 nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X12 G.t0 a_n10785_13139# VSS.t1 VSS.t0 nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X13 a_n12633_13089# a_n12405_13139# a_n12069_13139# VSS.t16 nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X14 a_n11457_13139# A.t1 E.t2 VSS.t13 nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X15 VSS.t3 B.t4 a_n11097_13463# VSS.t2 nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X16 E.t1 A.t2 a_n11709_13531# VDD.t13 pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X17 a_n11709_13531# a_n12405_13139# VDD.t19 VDD.t18 pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X18 a_n12405_13139# A.t3 VDD.t12 VDD.t11 pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X19 VDD.t17 a_n12405_13139# a_n12633_13089# VDD.t16 pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X20 VSS.t12 A.t4 a_n10617_13139# VSS.t11 nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X21 a_n12633_13089# B.t5 VDD.t3 VDD.t2 pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X22 G.t1 a_n10785_13139# VDD.t1 VDD.t0 pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X23 VDD.t15 A.t5 a_n10785_13139# VDD.t14 pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
R0 B.n0 B.t0 208.05
R1 B.t5 B.n0 177.391
R2 B.t3 B.t1 62.4155
R3 B.t0 B.t4 56.645
R4 B.n0 B.t3 35.0405
R5 B.n1 B.t5 30.0244
R6 B.n1 B.t2 21.7545
R7 B B.n1 12.5363
R8 VDD.n20 VDD.n5 337.079
R9 VDD.n22 VDD.t8 320.226
R10 VDD.n27 VDD.t14 286.517
R11 VDD.n11 VDD.t2 286.517
R12 VDD.t18 VDD.t13 235.956
R13 VDD.n21 VDD.t4 219.101
R14 VDD.n27 VDD.t6 185.393
R15 VDD.n26 VDD.t9 185.393
R16 VDD.t16 VDD.n15 185.393
R17 VDD.n11 VDD.t11 185.393
R18 VDD.t6 VDD.n3 154.617
R19 VDD.t11 VDD.n10 154.617
R20 VDD.n22 VDD.t9 151.685
R21 VDD.n16 VDD.t16 151.685
R22 VDD.t4 VDD.n20 117.978
R23 VDD.n16 VDD.t18 84.2702
R24 VDD.n3 VDD.t0 61.7474
R25 VDD.n10 VDD.t20 61.7474
R26 VDD.t14 VDD.n26 50.5623
R27 VDD.n15 VDD.t2 50.5623
R28 VDD.t8 VDD.n21 16.8544
R29 VDD.t13 VDD.n5 16.8544
R30 VDD.n28 VDD.n27 12.6005
R31 VDD.n26 VDD.n25 12.6005
R32 VDD.n23 VDD.n22 12.6005
R33 VDD.n21 VDD.n4 12.6005
R34 VDD.n20 VDD.n19 12.6005
R35 VDD.n18 VDD.n5 12.6005
R36 VDD.n17 VDD.n16 12.6005
R37 VDD.n15 VDD.n14 12.6005
R38 VDD.n12 VDD.n11 12.6005
R39 VDD.n3 VDD.n1 9.24875
R40 VDD.n10 VDD.n9 9.24875
R41 VDD.n19 VDD.t5 3.3856
R42 VDD.n13 VDD.t3 3.3856
R43 VDD.n24 VDD.t10 3.3856
R44 VDD.n2 VDD.t15 3.3856
R45 VDD.n9 VDD.n8 2.27383
R46 VDD.n7 VDD.n6 2.27383
R47 VDD.n1 VDD.n0 2.27383
R48 VDD.n8 VDD.t12 1.11226
R49 VDD.n8 VDD.t21 1.11226
R50 VDD.n6 VDD.t19 1.11226
R51 VDD.n6 VDD.t17 1.11226
R52 VDD.n0 VDD.t1 1.11226
R53 VDD.n0 VDD.t7 1.11226
R54 VDD.n23 VDD.n4 0.154786
R55 VDD.n19 VDD.n4 0.154786
R56 VDD.n19 VDD.n18 0.154786
R57 VDD.n18 VDD.n17 0.154786
R58 VDD.n25 VDD.n24 0.139357
R59 VDD.n14 VDD.n7 0.139357
R60 VDD.n12 VDD.n9 0.139357
R61 VDD.n28 VDD.n2 0.0776429
R62 VDD.n25 VDD.n2 0.0776429
R63 VDD.n14 VDD.n13 0.0776429
R64 VDD.n13 VDD.n12 0.0776429
R65 VDD VDD.n28 0.0744286
R66 VDD VDD.n1 0.0654286
R67 VDD.n24 VDD.n23 0.0159286
R68 VDD.n17 VDD.n7 0.0159286
R69 A.n0 A.t0 186.758
R70 A.t4 A.n0 186.758
R71 A.t1 A.t2 62.4155
R72 A.t0 A.t3 56.645
R73 A.n1 A.t5 30.0244
R74 A.n0 A.t1 24.6988
R75 A.n1 A.t4 21.7545
R76 A A.n1 12.5374
R77 VSS.n22 VSS.t10 1118.28
R78 VSS.n16 VSS.t16 1118.28
R79 VSS.n26 VSS.t11 1048.39
R80 VSS.t4 VSS.n12 1048.39
R81 VSS.n18 VSS.t6 978.495
R82 VSS.n18 VSS.t13 978.495
R83 VSS.n26 VSS.t2 908.602
R84 VSS.n12 VSS.t14 908.602
R85 VSS.n22 VSS.t8 838.711
R86 VSS.t17 VSS.n16 838.711
R87 VSS.t8 VSS.n21 559.14
R88 VSS.n17 VSS.t17 559.14
R89 VSS.t2 VSS.n3 492.834
R90 VSS.n9 VSS.t14 492.834
R91 VSS.n21 VSS.t6 419.356
R92 VSS.t13 VSS.n17 419.356
R93 VSS.t11 VSS.n25 349.462
R94 VSS.n13 VSS.t4 349.462
R95 VSS.n3 VSS.t0 316.954
R96 VSS.n9 VSS.t18 316.954
R97 VSS.n25 VSS.t10 279.57
R98 VSS.n13 VSS.t16 279.57
R99 VSS.n27 VSS.n26 10.4005
R100 VSS.n25 VSS.n24 10.4005
R101 VSS.n23 VSS.n22 10.4005
R102 VSS.n21 VSS.n20 10.4005
R103 VSS.n19 VSS.n18 10.4005
R104 VSS.n17 VSS.n6 10.4005
R105 VSS.n16 VSS.n15 10.4005
R106 VSS.n14 VSS.n13 10.4005
R107 VSS.n12 VSS.n11 10.4005
R108 VSS.n2 VSS.t12 8.64956
R109 VSS.n7 VSS.t5 8.64956
R110 VSS.n3 VSS.n1 6.73853
R111 VSS.n10 VSS.n9 6.73853
R112 VSS.n10 VSS.n8 6.64838
R113 VSS.n1 VSS.n0 6.64838
R114 VSS.n5 VSS.n4 6.64838
R115 VSS.n8 VSS.t15 2.00168
R116 VSS.n8 VSS.t19 2.00168
R117 VSS.n0 VSS.t1 2.00168
R118 VSS.n0 VSS.t3 2.00168
R119 VSS.n4 VSS.t9 2.00168
R120 VSS.n4 VSS.t7 2.00168
R121 VSS.n24 VSS.n23 0.154786
R122 VSS.n20 VSS.n19 0.154786
R123 VSS.n19 VSS.n6 0.154786
R124 VSS.n15 VSS.n6 0.154786
R125 VSS.n15 VSS.n14 0.154786
R126 VSS.n11 VSS.n10 0.154786
R127 VSS.n23 VSS.n5 0.147714
R128 VSS.n24 VSS.n2 0.0930714
R129 VSS.n14 VSS.n7 0.0930714
R130 VSS VSS.n1 0.0808571
R131 VSS VSS.n27 0.0744286
R132 VSS.n27 VSS.n2 0.0622143
R133 VSS.n11 VSS.n7 0.0622143
R134 VSS.n20 VSS.n5 0.00757143
R135 L.n0 L.t0 8.48448
R136 L L.n0 4.53959
R137 L.n0 L.t1 3.32871
R138 E E.n1 10.9908
R139 E.n0 E.t0 5.70523
R140 E.n0 E.t1 5.09613
R141 E.n1 E.t2 2.00168
R142 E.n1 E.t3 2.00168
R143 E E.n0 0.3485
R144 G.n0 G.t0 8.48457
R145 G G.n0 4.54595
R146 G.n0 G.t1 3.32566
C0 a_n11793_13139# a_n11709_13531# 0.01886f
C1 a_n11793_13139# a_n12405_13139# 0.05602f
C2 E a_n12633_13089# 0.02613f
C3 E a_n10785_13139# 0.01535f
C4 a_n11709_13531# a_n12633_13089# 0.0102f
C5 a_n12405_13139# a_n12633_13089# 0.46444f
C6 G VDD 0.22106f
C7 E a_n11097_13463# 0.05771f
C8 a_n11709_13531# a_n11097_13463# 0.02347f
C9 a_n11793_13139# B 0.01507f
C10 a_n11793_13139# a_n11457_13139# 0.20116f
C11 a_n12633_13089# VDD 0.44114f
C12 VDD a_n10785_13139# 0.44013f
C13 a_n12405_13139# L 0.01676f
C14 B a_n12633_13089# 0.17698f
C15 B a_n10785_13139# 0.05981f
C16 a_n11457_13139# a_n10785_13139# 0.11011f
C17 a_n11097_13463# VDD 0.66461f
C18 E a_n11709_13531# 0.59619f
C19 E a_n12405_13139# 0.06009f
C20 a_n11709_13531# a_n12405_13139# 0.02978f
C21 a_n11097_13463# B 0.11991f
C22 a_n11097_13463# a_n11457_13139# 0.09361f
C23 L VDD 0.22013f
C24 E VDD 0.56789f
C25 a_n11709_13531# VDD 0.44627f
C26 a_n12405_13139# VDD 0.6383f
C27 E B 0.0461f
C28 E a_n11457_13139# 0.12222f
C29 a_n11709_13531# B 0.04784f
C30 a_n11709_13531# a_n11457_13139# 0.30402f
C31 a_n12405_13139# B 0.24058f
C32 a_n11793_13139# A 0.03927f
C33 B VDD 1.58027f
C34 A a_n12633_13089# 0.0641f
C35 a_n11457_13139# VDD 0.02145f
C36 A a_n10785_13139# 0.18129f
C37 a_n11457_13139# B 0.02796f
C38 a_n11097_13463# A 0.24484f
C39 G a_n10785_13139# 0.20808f
C40 a_n11793_13139# a_n12633_13089# 0.10618f
C41 E A 0.05479f
C42 a_n11709_13531# A 0.04922f
C43 a_n12405_13139# A 0.12379f
C44 G a_n11097_13463# 0.01615f
C45 a_n11097_13463# a_n10785_13139# 0.49374f
C46 A VDD 0.42744f
C47 a_n12633_13089# L 0.20095f
C48 A B 0.1305f
C49 a_n11793_13139# E 0.19862f
C50 A a_n11457_13139# 0.01778f
C51 G VSS 0.29645f
C52 E VSS 0.22034f
C53 L VSS 0.30148f
C54 A VSS 1.92133f
C55 B VSS 0.82804f
C56 VDD VSS 7.18787f
C57 a_n11457_13139# VSS 0.24f
C58 a_n11793_13139# VSS 0.7516f
C59 a_n11709_13531# VSS 0.01037f
C60 a_n10785_13139# VSS 0.73563f
C61 a_n11097_13463# VSS 0.72346f
C62 a_n12405_13139# VSS 0.70755f
C63 a_n12633_13089# VSS 0.72971f
.ends

