magic
tech gf180mcuD
timestamp 1755250584
<< nwell >>
rect 0 63 253 127
rect 258 82 392 146
rect 0 -113 255 -49
rect 258 -50 322 14
<< nmos >>
rect 277 40 283 57
rect 294 40 300 57
rect 310 40 316 57
rect 333 40 339 57
rect 349 40 355 57
rect 366 40 372 57
rect 19 21 25 38
rect 36 21 42 38
rect 49 21 55 38
rect 72 21 78 38
rect 85 21 91 38
rect 102 21 108 38
rect 147 21 153 38
rect 164 21 170 38
rect 213 21 219 38
rect 224 21 230 38
rect 19 -24 25 -7
rect 36 -24 42 -7
rect 52 -24 58 -7
rect 75 -24 81 -7
rect 91 -24 97 -7
rect 108 -24 114 -7
rect 150 -24 156 -7
rect 161 -24 167 -7
rect 210 -24 216 -7
rect 227 -24 233 -7
rect 277 -92 283 -75
rect 294 -92 300 -75
<< pmos >>
rect 19 72 25 106
rect 36 72 42 106
rect 49 72 55 106
rect 72 72 78 106
rect 85 72 91 106
rect 102 72 108 106
rect 150 72 156 106
rect 161 72 167 106
rect 210 72 216 106
rect 227 72 233 106
rect 277 91 283 125
rect 294 91 300 125
rect 310 91 316 125
rect 333 91 339 125
rect 349 91 355 125
rect 366 91 372 125
rect 280 -41 286 -7
rect 291 -41 297 -7
rect 19 -92 25 -58
rect 36 -92 42 -58
rect 52 -92 58 -58
rect 75 -92 81 -58
rect 91 -92 97 -58
rect 108 -92 114 -58
rect 147 -92 153 -58
rect 164 -92 170 -58
rect 213 -92 219 -58
rect 224 -92 230 -58
<< ndiff >>
rect 58 38 68 39
rect 267 55 277 57
rect 267 42 269 55
rect 274 42 277 55
rect 267 40 277 42
rect 283 55 294 57
rect 283 42 286 55
rect 291 42 294 55
rect 283 40 294 42
rect 300 40 310 57
rect 316 47 333 57
rect 316 42 322 47
rect 327 42 333 47
rect 316 40 333 42
rect 339 40 349 57
rect 355 54 366 57
rect 355 42 358 54
rect 363 42 366 54
rect 355 40 366 42
rect 372 55 382 57
rect 372 42 375 55
rect 380 42 382 55
rect 372 40 382 42
rect 9 36 19 38
rect 9 23 11 36
rect 16 23 19 36
rect 9 21 19 23
rect 25 36 36 38
rect 25 23 28 36
rect 33 23 36 36
rect 25 21 36 23
rect 42 21 49 38
rect 55 37 72 38
rect 55 23 61 37
rect 66 23 72 37
rect 55 21 72 23
rect 78 21 85 38
rect 91 36 102 38
rect 91 23 94 36
rect 99 23 102 36
rect 91 21 102 23
rect 108 36 118 38
rect 108 23 111 36
rect 116 23 118 36
rect 108 21 118 23
rect 137 36 147 38
rect 137 23 139 36
rect 144 23 147 36
rect 137 21 147 23
rect 153 36 164 38
rect 153 23 156 36
rect 161 23 164 36
rect 153 21 164 23
rect 170 36 180 38
rect 170 23 173 36
rect 178 23 180 36
rect 170 21 180 23
rect 203 29 213 38
rect 203 23 205 29
rect 210 23 213 29
rect 203 21 213 23
rect 219 21 224 38
rect 230 36 240 38
rect 230 23 233 36
rect 238 23 240 36
rect 230 21 240 23
rect 9 -9 19 -7
rect 9 -22 11 -9
rect 16 -22 19 -9
rect 9 -24 19 -22
rect 25 -9 36 -7
rect 25 -22 28 -9
rect 33 -22 36 -9
rect 25 -24 36 -22
rect 42 -24 52 -7
rect 58 -9 75 -7
rect 58 -14 64 -9
rect 69 -14 75 -9
rect 58 -24 75 -14
rect 81 -24 91 -7
rect 97 -9 108 -7
rect 97 -21 100 -9
rect 105 -21 108 -9
rect 97 -24 108 -21
rect 114 -9 124 -7
rect 114 -22 117 -9
rect 122 -22 124 -9
rect 114 -24 124 -22
rect 140 -9 150 -7
rect 140 -15 142 -9
rect 147 -15 150 -9
rect 140 -24 150 -15
rect 156 -24 161 -7
rect 167 -9 177 -7
rect 167 -22 170 -9
rect 175 -22 177 -9
rect 167 -24 177 -22
rect 200 -9 210 -7
rect 200 -22 202 -9
rect 207 -22 210 -9
rect 200 -24 210 -22
rect 216 -9 227 -7
rect 216 -22 219 -9
rect 224 -22 227 -9
rect 216 -24 227 -22
rect 233 -9 243 -7
rect 233 -22 236 -9
rect 241 -22 243 -9
rect 233 -24 243 -22
rect 267 -77 277 -75
rect 267 -90 269 -77
rect 274 -90 277 -77
rect 267 -92 277 -90
rect 283 -77 294 -75
rect 283 -90 286 -77
rect 291 -90 294 -77
rect 283 -92 294 -90
rect 300 -77 310 -75
rect 300 -90 303 -77
rect 308 -90 310 -77
rect 300 -92 310 -90
<< pdiff >>
rect 267 123 277 125
rect 9 104 19 106
rect 9 96 11 104
rect 16 96 19 104
rect 9 72 19 96
rect 25 104 36 106
rect 25 96 28 104
rect 33 96 36 104
rect 25 72 36 96
rect 42 72 49 106
rect 55 104 72 106
rect 55 96 61 104
rect 66 96 72 104
rect 55 72 72 96
rect 78 72 85 106
rect 91 104 102 106
rect 91 96 94 104
rect 99 96 102 104
rect 91 72 102 96
rect 108 104 118 106
rect 108 96 111 104
rect 116 96 118 104
rect 108 72 118 96
rect 140 104 150 106
rect 140 74 142 104
rect 147 74 150 104
rect 140 72 150 74
rect 156 72 161 106
rect 167 104 177 106
rect 167 81 170 104
rect 175 81 177 104
rect 167 72 177 81
rect 200 104 210 106
rect 200 74 202 104
rect 207 74 210 104
rect 200 72 210 74
rect 216 104 227 106
rect 216 79 219 104
rect 224 79 227 104
rect 216 72 227 79
rect 233 104 243 106
rect 233 74 236 104
rect 241 74 243 104
rect 267 93 269 123
rect 274 93 277 123
rect 267 91 277 93
rect 283 123 294 125
rect 283 99 286 123
rect 291 99 294 123
rect 283 91 294 99
rect 300 91 310 125
rect 316 123 333 125
rect 316 118 322 123
rect 327 118 333 123
rect 316 91 333 118
rect 339 91 349 125
rect 355 123 366 125
rect 355 99 358 123
rect 363 99 366 123
rect 355 91 366 99
rect 372 123 382 125
rect 372 93 375 123
rect 380 93 382 123
rect 372 91 382 93
rect 233 72 243 74
rect 270 -9 280 -7
rect 270 -39 272 -9
rect 277 -39 280 -9
rect 270 -41 280 -39
rect 286 -41 291 -7
rect 297 -9 307 -7
rect 297 -32 300 -9
rect 305 -32 307 -9
rect 297 -41 307 -32
rect 9 -60 19 -58
rect 9 -90 11 -60
rect 16 -90 19 -60
rect 9 -92 19 -90
rect 25 -66 36 -58
rect 25 -90 28 -66
rect 33 -90 36 -66
rect 25 -92 36 -90
rect 42 -92 52 -58
rect 58 -85 75 -58
rect 58 -90 64 -85
rect 69 -90 75 -85
rect 58 -92 75 -90
rect 81 -92 91 -58
rect 97 -66 108 -58
rect 97 -90 100 -66
rect 105 -90 108 -66
rect 97 -92 108 -90
rect 114 -60 124 -58
rect 114 -90 117 -60
rect 122 -90 124 -60
rect 114 -92 124 -90
rect 137 -60 147 -58
rect 137 -90 139 -60
rect 144 -90 147 -60
rect 137 -92 147 -90
rect 153 -65 164 -58
rect 153 -90 156 -65
rect 161 -90 164 -65
rect 153 -92 164 -90
rect 170 -60 180 -58
rect 170 -90 173 -60
rect 178 -90 180 -60
rect 170 -92 180 -90
rect 203 -60 213 -58
rect 203 -90 205 -60
rect 210 -90 213 -60
rect 203 -92 213 -90
rect 219 -92 224 -58
rect 230 -67 240 -58
rect 230 -90 233 -67
rect 238 -90 240 -67
rect 230 -92 240 -90
<< ndiffc >>
rect 269 42 274 55
rect 286 42 291 55
rect 322 42 327 47
rect 358 42 363 54
rect 375 42 380 55
rect 11 23 16 36
rect 28 23 33 36
rect 61 23 66 37
rect 94 23 99 36
rect 111 23 116 36
rect 139 23 144 36
rect 156 23 161 36
rect 173 23 178 36
rect 205 23 210 29
rect 233 23 238 36
rect 11 -22 16 -9
rect 28 -22 33 -9
rect 64 -14 69 -9
rect 100 -21 105 -9
rect 117 -22 122 -9
rect 142 -15 147 -9
rect 170 -22 175 -9
rect 202 -22 207 -9
rect 219 -22 224 -9
rect 236 -22 241 -9
rect 269 -90 274 -77
rect 286 -90 291 -77
rect 303 -90 308 -77
<< pdiffc >>
rect 11 96 16 104
rect 28 96 33 104
rect 61 96 66 104
rect 94 96 99 104
rect 111 96 116 104
rect 142 74 147 104
rect 170 81 175 104
rect 202 74 207 104
rect 219 79 224 104
rect 236 74 241 104
rect 269 93 274 123
rect 286 99 291 123
rect 322 118 327 123
rect 358 99 363 123
rect 375 93 380 123
rect 272 -39 277 -9
rect 300 -32 305 -9
rect 11 -90 16 -60
rect 28 -90 33 -66
rect 64 -90 69 -85
rect 100 -90 105 -66
rect 117 -90 122 -60
rect 139 -90 144 -60
rect 156 -90 161 -65
rect 173 -90 178 -60
rect 205 -90 210 -60
rect 233 -90 238 -67
<< psubdiff >>
rect 264 31 279 33
rect 264 26 269 31
rect 274 26 279 31
rect 264 24 279 26
rect 288 31 303 33
rect 288 26 293 31
rect 298 26 303 31
rect 288 24 303 26
rect 312 31 327 33
rect 312 26 317 31
rect 322 26 327 31
rect 312 24 327 26
rect 336 31 351 33
rect 336 26 341 31
rect 346 26 351 31
rect 336 24 351 26
rect 360 31 375 33
rect 360 26 365 31
rect 370 26 375 31
rect 360 24 375 26
rect 6 12 21 14
rect 6 2 11 12
rect 16 2 21 12
rect 6 0 21 2
rect 30 12 45 14
rect 30 2 35 12
rect 40 2 45 12
rect 30 0 45 2
rect 54 12 69 14
rect 54 2 59 12
rect 64 2 69 12
rect 54 0 69 2
rect 78 12 93 14
rect 78 2 83 12
rect 88 2 93 12
rect 78 0 93 2
rect 102 12 117 14
rect 102 2 107 12
rect 112 2 117 12
rect 102 0 117 2
rect 134 12 149 14
rect 134 2 139 12
rect 144 2 149 12
rect 134 0 149 2
rect 158 12 173 14
rect 158 2 163 12
rect 168 2 173 12
rect 158 0 173 2
rect 197 12 212 14
rect 197 2 202 12
rect 207 2 212 12
rect 197 0 212 2
rect 221 12 236 14
rect 221 2 226 12
rect 231 2 236 12
rect 221 0 236 2
rect 264 -101 279 -99
rect 264 -106 269 -101
rect 274 -106 279 -101
rect 264 -108 279 -106
rect 288 -101 303 -99
rect 288 -106 293 -101
rect 298 -106 303 -101
rect 288 -108 303 -106
<< nsubdiff >>
rect 264 139 279 141
rect 264 134 269 139
rect 274 134 279 139
rect 264 132 279 134
rect 288 139 303 141
rect 288 134 293 139
rect 298 134 303 139
rect 288 132 303 134
rect 312 139 327 141
rect 312 134 317 139
rect 322 134 327 139
rect 312 132 327 134
rect 336 139 351 141
rect 336 134 341 139
rect 346 134 351 139
rect 336 132 351 134
rect 360 139 375 141
rect 360 134 365 139
rect 370 134 375 139
rect 360 132 375 134
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
rect 54 120 69 122
rect 54 115 59 120
rect 64 115 69 120
rect 54 113 69 115
rect 78 120 93 122
rect 78 115 83 120
rect 88 115 93 120
rect 78 113 93 115
rect 102 120 117 122
rect 102 115 107 120
rect 112 115 117 120
rect 102 113 117 115
rect 134 120 149 122
rect 134 115 139 120
rect 144 115 149 120
rect 134 113 149 115
rect 158 120 173 122
rect 158 115 163 120
rect 168 115 173 120
rect 158 113 173 115
rect 197 120 212 122
rect 197 115 202 120
rect 207 115 212 120
rect 197 113 212 115
rect 221 120 236 122
rect 221 115 226 120
rect 231 115 236 120
rect 221 113 236 115
rect 264 7 279 9
rect 264 2 269 7
rect 274 2 279 7
rect 264 0 279 2
rect 288 7 303 9
rect 288 2 293 7
rect 298 2 303 7
rect 288 0 303 2
rect 6 -101 21 -99
rect 6 -106 11 -101
rect 16 -106 21 -101
rect 6 -108 21 -106
rect 30 -101 45 -99
rect 30 -106 35 -101
rect 40 -106 45 -101
rect 30 -108 45 -106
rect 54 -101 69 -99
rect 54 -106 59 -101
rect 64 -106 69 -101
rect 54 -108 69 -106
rect 78 -101 93 -99
rect 78 -106 83 -101
rect 88 -106 93 -101
rect 78 -108 93 -106
rect 102 -101 117 -99
rect 102 -106 107 -101
rect 112 -106 117 -101
rect 102 -108 117 -106
rect 134 -101 149 -99
rect 134 -106 139 -101
rect 144 -106 149 -101
rect 134 -108 149 -106
rect 158 -101 173 -99
rect 158 -106 163 -101
rect 168 -106 173 -101
rect 158 -108 173 -106
rect 197 -101 212 -99
rect 197 -106 202 -101
rect 207 -106 212 -101
rect 197 -108 212 -106
rect 221 -101 236 -99
rect 221 -106 226 -101
rect 231 -106 236 -101
rect 221 -108 236 -106
<< psubdiffcont >>
rect 269 26 274 31
rect 293 26 298 31
rect 317 26 322 31
rect 341 26 346 31
rect 365 26 370 31
rect 11 2 16 12
rect 35 2 40 12
rect 59 2 64 12
rect 83 2 88 12
rect 107 2 112 12
rect 139 2 144 12
rect 163 2 168 12
rect 202 2 207 12
rect 226 2 231 12
rect 269 -106 274 -101
rect 293 -106 298 -101
<< nsubdiffcont >>
rect 269 134 274 139
rect 293 134 298 139
rect 317 134 322 139
rect 341 134 346 139
rect 365 134 370 139
rect 11 115 16 120
rect 35 115 40 120
rect 59 115 64 120
rect 83 115 88 120
rect 107 115 112 120
rect 139 115 144 120
rect 163 115 168 120
rect 202 115 207 120
rect 226 115 231 120
rect 269 2 274 7
rect 293 2 298 7
rect 11 -106 16 -101
rect 35 -106 40 -101
rect 59 -106 64 -101
rect 83 -106 88 -101
rect 107 -106 112 -101
rect 139 -106 144 -101
rect 163 -106 168 -101
rect 202 -106 207 -101
rect 226 -106 231 -101
<< polysilicon >>
rect 277 125 283 130
rect 294 125 300 130
rect 310 125 316 130
rect 333 125 339 130
rect 349 125 355 130
rect 366 125 372 130
rect 19 106 25 111
rect 36 106 42 111
rect 49 106 55 111
rect 72 106 78 111
rect 85 106 91 111
rect 102 106 108 111
rect 150 106 156 111
rect 161 106 167 111
rect 210 106 216 111
rect 227 106 233 111
rect 277 89 283 91
rect 294 89 300 91
rect 277 84 300 89
rect 310 89 316 91
rect 333 89 339 91
rect 310 87 320 89
rect 277 73 283 84
rect 310 82 312 87
rect 318 82 320 87
rect 310 80 320 82
rect 329 87 339 89
rect 329 81 331 87
rect 337 81 339 87
rect 349 89 355 91
rect 366 89 372 91
rect 349 84 372 89
rect 329 79 339 81
rect 19 54 25 72
rect 36 70 42 72
rect 31 68 42 70
rect 31 62 33 68
rect 39 62 42 68
rect 31 60 42 62
rect 49 70 55 72
rect 72 70 78 72
rect 85 70 91 72
rect 102 70 108 72
rect 49 68 63 70
rect 49 62 55 68
rect 61 62 63 68
rect 49 60 63 62
rect 70 68 80 70
rect 70 62 72 68
rect 78 62 80 68
rect 85 65 108 70
rect 150 68 156 72
rect 70 60 80 62
rect 19 52 35 54
rect 19 46 27 52
rect 33 51 35 52
rect 33 46 42 51
rect 19 44 42 46
rect 19 38 25 44
rect 36 38 42 44
rect 49 38 55 60
rect 102 54 108 65
rect 147 63 156 68
rect 161 69 167 72
rect 161 67 170 69
rect 161 65 178 67
rect 161 63 170 65
rect 147 54 153 63
rect 60 52 70 54
rect 91 52 108 54
rect 60 46 62 52
rect 68 46 78 52
rect 91 49 93 52
rect 60 44 78 46
rect 72 38 78 44
rect 85 46 93 49
rect 99 46 108 52
rect 85 44 108 46
rect 139 52 153 54
rect 139 46 142 52
rect 148 46 153 52
rect 139 44 153 46
rect 85 38 91 44
rect 102 38 108 44
rect 147 38 153 44
rect 164 59 170 63
rect 176 59 178 65
rect 164 57 178 59
rect 164 38 170 57
rect 210 54 216 72
rect 202 52 216 54
rect 202 46 205 52
rect 211 46 216 52
rect 202 44 216 46
rect 210 43 216 44
rect 227 67 233 72
rect 277 71 290 73
rect 227 65 241 67
rect 227 59 233 65
rect 239 59 241 65
rect 227 57 241 59
rect 277 65 282 71
rect 288 65 290 71
rect 277 63 290 65
rect 305 67 316 69
rect 277 59 300 63
rect 305 61 307 67
rect 313 61 316 67
rect 305 59 316 61
rect 277 57 283 59
rect 294 57 300 59
rect 310 57 316 59
rect 333 57 339 79
rect 345 77 355 79
rect 345 72 347 77
rect 353 72 355 77
rect 366 73 372 84
rect 345 70 355 72
rect 349 57 355 70
rect 360 71 372 73
rect 360 65 362 71
rect 368 65 372 71
rect 360 63 372 65
rect 366 57 372 63
rect 227 43 233 57
rect 210 40 219 43
rect 213 38 219 40
rect 224 40 233 43
rect 224 38 230 40
rect 277 35 283 40
rect 294 35 300 40
rect 310 35 316 40
rect 333 35 339 40
rect 349 35 355 40
rect 366 35 372 40
rect 19 16 25 21
rect 36 16 42 21
rect 49 16 55 21
rect 72 16 78 21
rect 85 16 91 21
rect 102 16 108 21
rect 147 16 153 21
rect 164 16 170 21
rect 213 16 219 21
rect 224 16 230 21
rect 19 -7 25 -2
rect 36 -7 42 -2
rect 52 -7 58 -2
rect 75 -7 81 -2
rect 91 -7 97 -2
rect 108 -7 114 -2
rect 150 -7 156 -2
rect 161 -7 167 -2
rect 210 -7 216 -2
rect 227 -7 233 -2
rect 280 -7 286 -2
rect 291 -7 297 -2
rect 19 -26 25 -24
rect 36 -26 42 -24
rect 52 -26 58 -24
rect 19 -30 42 -26
rect 47 -28 58 -26
rect 19 -32 32 -30
rect 19 -38 24 -32
rect 30 -38 32 -32
rect 47 -34 49 -28
rect 55 -34 58 -28
rect 47 -36 58 -34
rect 19 -40 32 -38
rect 19 -51 25 -40
rect 75 -46 81 -24
rect 91 -37 97 -24
rect 108 -30 114 -24
rect 150 -26 156 -24
rect 147 -29 156 -26
rect 161 -26 167 -24
rect 161 -29 170 -26
rect 147 -30 153 -29
rect 87 -39 97 -37
rect 87 -44 89 -39
rect 95 -44 97 -39
rect 102 -32 114 -30
rect 102 -38 104 -32
rect 110 -38 114 -32
rect 102 -40 114 -38
rect 139 -32 153 -30
rect 139 -38 142 -32
rect 148 -38 153 -32
rect 139 -40 153 -38
rect 87 -46 97 -44
rect 52 -49 62 -47
rect 19 -56 42 -51
rect 19 -58 25 -56
rect 36 -58 42 -56
rect 52 -54 54 -49
rect 60 -54 62 -49
rect 52 -56 62 -54
rect 71 -48 81 -46
rect 71 -54 73 -48
rect 79 -54 81 -48
rect 108 -51 114 -40
rect 71 -56 81 -54
rect 52 -58 58 -56
rect 75 -58 81 -56
rect 91 -56 114 -51
rect 91 -58 97 -56
rect 108 -58 114 -56
rect 147 -58 153 -40
rect 164 -43 170 -29
rect 210 -30 216 -24
rect 202 -32 216 -30
rect 202 -38 205 -32
rect 211 -38 216 -32
rect 202 -40 216 -38
rect 164 -45 178 -43
rect 164 -51 170 -45
rect 176 -51 178 -45
rect 164 -53 178 -51
rect 210 -49 216 -40
rect 227 -43 233 -24
rect 227 -45 241 -43
rect 280 -45 286 -41
rect 227 -49 233 -45
rect 164 -58 170 -53
rect 210 -54 219 -49
rect 213 -58 219 -54
rect 224 -51 233 -49
rect 239 -51 241 -45
rect 224 -53 241 -51
rect 277 -50 286 -45
rect 291 -44 297 -41
rect 291 -46 300 -44
rect 291 -48 308 -46
rect 291 -50 300 -48
rect 224 -55 233 -53
rect 224 -58 230 -55
rect 277 -59 283 -50
rect 269 -61 283 -59
rect 269 -67 272 -61
rect 278 -67 283 -61
rect 269 -69 283 -67
rect 277 -75 283 -69
rect 294 -54 300 -50
rect 306 -54 308 -48
rect 294 -56 308 -54
rect 294 -75 300 -56
rect 19 -97 25 -92
rect 36 -97 42 -92
rect 52 -97 58 -92
rect 75 -97 81 -92
rect 91 -97 97 -92
rect 108 -97 114 -92
rect 147 -97 153 -92
rect 164 -97 170 -92
rect 213 -97 219 -92
rect 224 -97 230 -92
rect 277 -97 283 -92
rect 294 -97 300 -92
<< polycontact >>
rect 312 82 318 87
rect 331 81 337 87
rect 33 62 39 68
rect 55 62 61 68
rect 72 62 78 68
rect 27 46 33 52
rect 62 46 68 52
rect 93 46 99 52
rect 142 46 148 52
rect 170 59 176 65
rect 205 46 211 52
rect 233 59 239 65
rect 282 65 288 71
rect 307 61 313 67
rect 347 72 353 77
rect 362 65 368 71
rect 24 -38 30 -32
rect 49 -34 55 -28
rect 89 -44 95 -39
rect 104 -38 110 -32
rect 142 -38 148 -32
rect 54 -54 60 -49
rect 73 -54 79 -48
rect 205 -38 211 -32
rect 170 -51 176 -45
rect 233 -51 239 -45
rect 272 -67 278 -61
rect 300 -54 306 -48
<< metal1 >>
rect 258 139 392 146
rect 258 134 269 139
rect 274 134 293 139
rect 298 134 317 139
rect 322 134 341 139
rect 346 134 365 139
rect 370 134 392 139
rect 258 132 392 134
rect 0 120 253 127
rect 0 115 11 120
rect 16 115 35 120
rect 40 115 59 120
rect 64 115 83 120
rect 88 115 107 120
rect 112 115 139 120
rect 144 115 163 120
rect 168 115 202 120
rect 207 115 226 120
rect 231 115 253 120
rect 0 113 253 115
rect 269 123 274 125
rect 11 104 16 106
rect 11 68 16 96
rect 28 104 33 113
rect 61 104 66 106
rect 28 94 33 96
rect 60 96 61 97
rect 60 91 66 96
rect 94 104 99 113
rect 94 94 99 96
rect 111 104 116 106
rect 60 83 66 85
rect 111 78 116 96
rect 55 73 116 78
rect 55 68 61 73
rect 11 62 33 68
rect 39 62 48 68
rect 11 36 16 62
rect 42 52 48 62
rect 70 62 72 68
rect 78 62 80 68
rect 55 60 61 62
rect 25 46 27 52
rect 33 46 35 52
rect 42 46 62 52
rect 68 46 70 52
rect 91 46 93 52
rect 99 46 101 52
rect 60 39 66 41
rect 11 21 16 23
rect 28 36 33 38
rect 60 30 61 33
rect 28 14 33 23
rect 61 21 66 23
rect 94 36 99 38
rect 94 14 99 23
rect 111 36 116 73
rect 142 104 147 113
rect 170 104 175 106
rect 170 79 175 81
rect 156 78 175 79
rect 142 72 147 74
rect 154 72 156 78
rect 162 74 175 78
rect 202 104 207 113
rect 219 104 224 106
rect 219 78 224 79
rect 236 104 241 113
rect 162 72 164 74
rect 202 72 207 74
rect 217 72 219 78
rect 225 72 227 78
rect 236 72 241 74
rect 286 123 291 132
rect 322 123 327 125
rect 322 112 327 118
rect 321 110 327 112
rect 358 123 363 132
rect 319 104 321 110
rect 327 104 329 110
rect 286 97 291 99
rect 269 86 274 93
rect 312 94 352 99
rect 358 97 363 99
rect 375 123 380 125
rect 312 87 318 94
rect 347 89 352 94
rect 375 89 380 93
rect 331 87 337 89
rect 269 81 305 86
rect 310 82 312 87
rect 318 82 320 87
rect 140 46 142 52
rect 148 46 150 52
rect 111 21 116 23
rect 139 36 144 38
rect 139 14 144 23
rect 156 36 161 72
rect 168 59 170 65
rect 176 59 178 65
rect 203 46 205 52
rect 211 46 213 52
rect 156 21 161 23
rect 173 36 178 38
rect 219 37 224 72
rect 231 59 233 65
rect 239 59 241 65
rect 269 55 274 81
rect 299 77 305 81
rect 331 77 337 81
rect 347 83 380 89
rect 347 78 353 83
rect 299 72 337 77
rect 345 77 355 78
rect 345 72 347 77
rect 353 72 355 77
rect 280 65 282 71
rect 288 65 290 71
rect 360 67 362 71
rect 305 61 307 67
rect 313 65 362 67
rect 368 65 370 71
rect 313 61 367 65
rect 269 40 274 42
rect 286 55 291 57
rect 321 55 327 56
rect 319 49 321 55
rect 327 49 329 55
rect 358 54 363 56
rect 321 47 327 49
rect 173 14 178 23
rect 205 32 224 37
rect 233 36 238 38
rect 205 29 210 32
rect 205 21 210 23
rect 286 33 291 42
rect 322 40 327 42
rect 358 33 363 42
rect 375 55 380 83
rect 375 40 380 42
rect 233 14 238 23
rect 258 31 392 33
rect 258 26 269 31
rect 274 26 293 31
rect 298 26 317 31
rect 322 26 341 31
rect 346 26 365 31
rect 370 26 392 31
rect 258 19 392 26
rect 0 12 255 14
rect 0 2 11 12
rect 16 2 35 12
rect 40 2 59 12
rect 64 2 83 12
rect 88 2 107 12
rect 112 2 139 12
rect 144 2 163 12
rect 168 2 202 12
rect 207 2 226 12
rect 231 2 255 12
rect 0 0 255 2
rect 258 7 322 14
rect 258 2 269 7
rect 274 2 293 7
rect 298 2 322 7
rect 258 0 322 2
rect 11 -9 16 -7
rect 11 -48 16 -22
rect 28 -9 33 0
rect 64 -9 69 -7
rect 63 -16 69 -14
rect 100 -9 105 0
rect 61 -22 63 -16
rect 69 -22 71 -16
rect 28 -24 33 -22
rect 63 -23 69 -22
rect 100 -23 105 -21
rect 117 -9 122 -7
rect 22 -38 24 -32
rect 30 -38 32 -32
rect 47 -34 49 -28
rect 55 -32 109 -28
rect 55 -34 104 -32
rect 102 -38 104 -34
rect 110 -38 112 -32
rect 41 -44 79 -39
rect 41 -48 47 -44
rect 11 -53 47 -48
rect 73 -48 79 -44
rect 87 -44 89 -39
rect 95 -44 97 -39
rect 87 -45 97 -44
rect 11 -60 16 -53
rect 52 -54 54 -49
rect 60 -54 62 -49
rect 54 -61 60 -54
rect 73 -56 79 -54
rect 89 -50 95 -45
rect 117 -50 122 -22
rect 142 -9 147 -7
rect 142 -18 147 -15
rect 170 -9 175 0
rect 142 -23 161 -18
rect 140 -38 142 -32
rect 148 -38 150 -32
rect 89 -56 122 -50
rect 89 -61 94 -56
rect 11 -92 16 -90
rect 28 -66 33 -64
rect 54 -66 94 -61
rect 117 -60 122 -56
rect 156 -58 161 -23
rect 170 -24 175 -22
rect 202 -9 207 0
rect 202 -24 207 -22
rect 219 -9 224 -7
rect 203 -38 205 -32
rect 211 -38 213 -32
rect 168 -51 170 -45
rect 176 -51 178 -45
rect 219 -58 224 -22
rect 236 -9 241 0
rect 236 -24 241 -22
rect 272 -9 277 0
rect 300 -9 305 -7
rect 300 -34 305 -32
rect 286 -35 305 -34
rect 272 -41 277 -39
rect 284 -41 286 -35
rect 292 -39 305 -35
rect 292 -41 294 -39
rect 231 -51 233 -45
rect 239 -51 241 -45
rect 100 -66 105 -64
rect 61 -77 63 -71
rect 69 -77 71 -71
rect 63 -79 69 -77
rect 28 -99 33 -90
rect 64 -85 69 -79
rect 64 -92 69 -90
rect 100 -99 105 -90
rect 117 -92 122 -90
rect 139 -60 144 -58
rect 154 -64 156 -58
rect 162 -64 164 -58
rect 173 -60 178 -58
rect 139 -99 144 -90
rect 156 -65 161 -64
rect 156 -92 161 -90
rect 173 -99 178 -90
rect 205 -60 210 -58
rect 217 -64 219 -58
rect 225 -60 227 -58
rect 225 -64 238 -60
rect 219 -65 238 -64
rect 205 -99 210 -90
rect 233 -67 238 -65
rect 270 -67 272 -61
rect 278 -67 280 -61
rect 233 -92 238 -90
rect 269 -77 274 -75
rect 269 -99 274 -90
rect 286 -77 291 -41
rect 298 -54 300 -48
rect 306 -54 308 -48
rect 286 -92 291 -90
rect 303 -77 308 -75
rect 303 -99 308 -90
rect 0 -101 255 -99
rect 0 -106 11 -101
rect 16 -106 35 -101
rect 40 -106 59 -101
rect 64 -106 83 -101
rect 88 -106 107 -101
rect 112 -106 139 -101
rect 144 -106 163 -101
rect 168 -106 202 -101
rect 207 -106 226 -101
rect 231 -106 255 -101
rect 0 -113 255 -106
rect 258 -101 322 -99
rect 258 -106 269 -101
rect 274 -106 293 -101
rect 298 -106 322 -101
rect 258 -113 322 -106
<< via1 >>
rect 60 85 66 91
rect 72 62 78 68
rect 27 46 33 52
rect 93 46 99 52
rect 60 37 66 39
rect 60 33 61 37
rect 61 33 66 37
rect 156 72 162 78
rect 219 72 225 78
rect 321 104 327 110
rect 142 46 148 52
rect 170 59 176 65
rect 205 46 211 52
rect 233 59 239 65
rect 282 65 288 71
rect 362 65 368 71
rect 321 49 327 55
rect 63 -22 69 -16
rect 24 -38 30 -32
rect 104 -38 110 -32
rect 142 -38 148 -32
rect 205 -38 211 -32
rect 170 -51 176 -45
rect 286 -41 292 -35
rect 233 -51 239 -45
rect 63 -77 69 -71
rect 156 -64 162 -58
rect 219 -64 225 -58
rect 272 -67 278 -61
rect 300 -54 306 -48
<< metal2 >>
rect 321 111 327 112
rect 320 110 328 111
rect 320 104 321 110
rect 327 104 328 110
rect 320 103 328 104
rect 60 92 66 97
rect 59 91 67 92
rect 59 85 60 91
rect 66 85 67 91
rect 59 84 67 85
rect 59 83 66 84
rect 27 53 33 54
rect 26 52 34 53
rect 26 46 27 52
rect 33 46 34 52
rect 26 45 34 46
rect 27 26 33 45
rect 59 40 65 83
rect 154 78 164 79
rect 154 72 156 78
rect 162 72 164 78
rect 154 71 164 72
rect 217 78 227 79
rect 217 72 219 78
rect 225 72 227 78
rect 217 71 227 72
rect 281 71 289 72
rect 72 69 79 70
rect 71 68 80 69
rect 71 62 72 68
rect 78 62 80 68
rect 71 61 80 62
rect 72 60 80 61
rect 58 39 68 40
rect 58 33 60 39
rect 66 33 68 39
rect 58 32 68 33
rect 74 26 80 60
rect 168 65 178 66
rect 168 59 170 65
rect 176 59 178 65
rect 168 58 178 59
rect 231 65 241 66
rect 280 65 282 71
rect 288 65 290 71
rect 231 59 233 65
rect 239 59 241 65
rect 281 64 289 65
rect 231 58 241 59
rect 321 56 327 103
rect 361 71 369 72
rect 360 65 362 71
rect 368 65 370 71
rect 361 64 369 65
rect 319 55 329 56
rect 93 53 99 54
rect 92 52 100 53
rect 140 52 150 53
rect 91 46 93 52
rect 99 46 101 52
rect 140 46 142 52
rect 148 46 150 52
rect 92 45 100 46
rect 140 45 150 46
rect 203 52 213 53
rect 203 46 205 52
rect 211 46 213 52
rect 319 49 321 55
rect 327 49 329 55
rect 319 48 329 49
rect 203 45 213 46
rect 93 44 99 45
rect 27 20 80 26
rect 61 -16 71 -15
rect 61 -22 63 -16
rect 69 -22 71 -16
rect 61 -23 71 -22
rect 23 -32 31 -31
rect 22 -38 24 -32
rect 30 -38 32 -32
rect 23 -39 31 -38
rect 63 -70 69 -23
rect 103 -32 111 -31
rect 140 -32 150 -31
rect 102 -38 104 -32
rect 110 -38 112 -32
rect 140 -38 142 -32
rect 148 -38 150 -32
rect 103 -39 111 -38
rect 140 -39 150 -38
rect 203 -32 213 -31
rect 203 -38 205 -32
rect 211 -38 213 -32
rect 203 -39 213 -38
rect 284 -35 294 -34
rect 284 -41 286 -35
rect 292 -41 294 -35
rect 284 -42 294 -41
rect 168 -45 178 -44
rect 168 -51 170 -45
rect 176 -51 178 -45
rect 168 -52 178 -51
rect 231 -45 241 -44
rect 231 -51 233 -45
rect 239 -51 241 -45
rect 231 -52 241 -51
rect 298 -48 308 -47
rect 298 -54 300 -48
rect 306 -54 308 -48
rect 298 -55 308 -54
rect 154 -58 164 -57
rect 154 -64 156 -58
rect 162 -64 164 -58
rect 154 -65 164 -64
rect 217 -58 227 -57
rect 217 -64 219 -58
rect 225 -64 227 -58
rect 217 -65 227 -64
rect 270 -61 280 -60
rect 270 -67 272 -61
rect 278 -67 280 -61
rect 270 -68 280 -67
rect 62 -71 70 -70
rect 62 -77 63 -71
rect 69 -77 70 -71
rect 62 -78 70 -77
rect 63 -79 69 -78
<< labels >>
rlabel metal2 30 49 30 49 1 my_nxor_0.A
rlabel metal2 63 87 63 87 1 my_nxor_0.Y
rlabel metal1 13 117 13 117 1 my_nxor_0.VDD
rlabel psubdiffcont 13 9 13 9 1 my_nxor_0.VSS
rlabel via1 27 -35 27 -35 5 my_xor_0.A
rlabel via1 107 -35 107 -35 5 my_xor_0.B
rlabel via1 66 -73 66 -73 5 my_xor_0.Y
rlabel nsubdiffcont 13 -104 13 -104 5 my_xor_0.VDD
rlabel psubdiffcont 13 4 13 4 5 my_xor_0.VSS
rlabel via1 145 -35 145 -35 5 my_nand_0.A
rlabel via1 173 -48 173 -48 5 my_nand_0.B
rlabel via1 159 -61 159 -61 5 my_nand_0.Y
rlabel nsubdiffcont 141 -104 141 -104 5 my_nand_0.VDD
rlabel psubdiffcont 141 5 141 5 5 my_nand_0.VSS
rlabel psubdiffcont 141 9 141 9 1 my_nor_0.VSS
rlabel nsubdiffcont 141 117 141 117 1 my_nor_0.VDD
rlabel via1 159 75 159 75 1 my_nor_0.Y
rlabel via1 173 62 173 62 1 my_nor_0.B
rlabel via1 145 49 145 49 1 my_nor_0.A
rlabel metal2 96 49 96 49 1 my_nxor_0.B
rlabel via1 208 -35 208 -35 5 my_nor_0.A
rlabel via1 236 -48 236 -48 5 my_nor_0.B
rlabel via1 222 -61 222 -61 5 my_nor_0.Y
rlabel nsubdiffcont 204 -103 204 -103 5 my_nor_0.VDD
rlabel psubdiffcont 204 5 204 5 5 my_nor_0.VSS
rlabel psubdiffcont 204 9 204 9 1 my_nand_0.VSS
rlabel nsubdiffcont 204 118 204 118 1 my_nand_0.VDD
rlabel via1 222 75 222 75 1 my_nand_0.Y
rlabel via1 236 62 236 62 1 my_nand_0.B
rlabel via1 208 49 208 49 1 my_nand_0.A
rlabel metal2 275 -64 275 -64 1 my_nor_0.A
rlabel metal2 303 -51 303 -51 1 my_nor_0.B
rlabel metal2 289 -38 289 -38 1 my_nor_0.Y
rlabel metal1 271 4 271 4 1 my_nor_0.VDD
rlabel metal1 271 -104 271 -104 1 my_nor_0.VSS
rlabel metal2 285 68 285 68 1 my_xor_0.A
rlabel metal2 365 68 365 68 1 my_xor_0.B
rlabel metal2 324 106 324 106 1 my_xor_0.Y
rlabel metal1 271 137 271 137 1 my_xor_0.VDD
rlabel metal1 271 29 271 29 1 my_xor_0.VSS
<< end >>
