* NGSPICE file created from gf180mcu_gp9t3v3__comp2_1.ext - technology: gf180mcuD

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

.subckt gf180mcu_gp9t3v3__comp2_1 L E G VDD VSS A B
X0 VDD B a_n11097_13463# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X1 a_n12405_13139# A VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X2 VSS B a_n11793_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X3 a_n10617_13139# a_n11097_13463# a_n10785_13139# VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X4 a_n10785_13139# a_n11097_13463# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X5 a_n12069_13139# B VSS VSS nfet_03v3 ad=0.102p pd=1.09u as=0.459p ps=2.78u w=0.85u l=0.3u
X6 VDD a_n12633_13089# L VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X7 E a_n11097_13463# a_n11709_13531# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X8 VSS a_n12633_13089# L VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X9 a_n11457_13139# a_n11097_13463# VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X10 a_n11709_13531# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X11 E a_n12405_13139# a_n11793_13139# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X12 G a_n10785_13139# VSS VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X13 a_n12633_13089# a_n12405_13139# a_n12069_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X14 a_n11457_13139# A E VSS nfet_03v3 ad=0.459p pd=2.78u as=0.2295p ps=1.39u w=0.85u l=0.3u
X15 VSS B a_n11097_13463# VSS nfet_03v3 ad=0.2295p pd=1.39u as=0.459p ps=2.78u w=0.85u l=0.3u
X16 E A a_n11709_13531# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X17 a_n11709_13531# a_n12405_13139# VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X18 a_n12405_13139# A VDD VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X19 VDD a_n12405_13139# a_n12633_13089# VDD pfet_03v3 ad=0.459p pd=2.24u as=0.459p ps=2.24u w=1.7u l=0.3u
X20 VSS A a_n10617_13139# VSS nfet_03v3 ad=0.459p pd=2.78u as=0.102p ps=1.09u w=0.85u l=0.3u
X21 a_n12633_13089# B VDD VDD pfet_03v3 ad=0.459p pd=2.24u as=0.918p ps=4.48u w=1.7u l=0.3u
X22 G a_n10785_13139# VDD VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
X23 VDD A a_n10785_13139# VDD pfet_03v3 ad=0.918p pd=4.48u as=0.459p ps=2.24u w=1.7u l=0.3u
.ends

