  X � 	   ) -� 	   ) - LIB  >A�7KƧ�9D�/��ZT � 	   ) -� 	   ) - gf180mcu_gp9t3v3__comp2_1         ,��!� G��!� ���*� ���*� G��!� G          ,��+� G��+� ���4c ���4c G��+� G          ,��w G��w ��� � ��� � G��w G          ,��5� G��5� ���>; ���>; G��5� G          ,��#�  ���#� ���,/ ���,/  ���#�  �          ,��-[  ���-[ ���4� ���4�  ���-[  �          ,��6  ���6 ���>� ���>�  ���6  �          ,���  ���� ���"W ���"W  ����  �          ,���  ���� ��� ���  ����  �          ,��� G��� ���K ���K G��� G          ,��'  ���' ���� ����  ���'  �          ,��!v )��!v ���$d ���$d )��!v )          ,��� )��� ���� ���� )��� )          ,�� )�� ��� ��� )�� )          ,��f )��f ���T ���T )��f )          ,��� )��� ���� ���� )��� )          ,��
 )��
 ���� ���� )��
 )          ,��8� )��8� ���;� ���;� )��8� )          ,��46 )��46 ���7$ ���7$ )��46 )          ,��/� )��/� ���2t ���2t )��/� )          ,��*� )��*� ���-� ���-� )��*� )          ,��&& )��&& ���) ���) )��&& )          ,��!v  ����!v  �a��$d  �a��$d  ����!v  ��          ,���  �����  �a���  �a���  �����  ��          ,��  ����  �a��  �a��  ����  ��          ,��f  ����f  �a��T  �a��T  ����f  ��          ,���  �����  �a���  �a���  �����  ��          ,��
  ����
  �a���  �a���  ����
  ��          ,��8�  ����8�  �a��;�  �a��;�  ����8�  ��          ,��46  ����46  �a��7$  �a��7$  ����46  ��          ,��/�  ����/�  �a��2t  �a��2t  ����/�  ��          ,��*�  ����*�  �a��-�  �a��-�  ����*�  ��          ,��&&  ����&&  �a��)  �a��)  ����&&  ��          ,��k ���k ���� ���� ���k �          ,��1 ���1 ���2G ���2G ���1 �          ,��:� ���:� ���< ���< ���:� �          ,��8#  ����8# }��9O }��9O  ����8#  ��          ,��1�  ����1� ���2� ���2�  ����1�  ��          ,��/w  ����/w }��0� }��0�  ����/w  ��          ,��;k  ����;k ���<� ���<�  ����;k  ��          ,��%�  ����%� }��&� }��&�  ����%�  ��          ,��(�  ����(� }��* }��*  ����(�  ��          ,���  ����� }��� }���  �����  ��          ,��  ���� ��� ; ��� ;  ����  ��          ,��	C  ����	C ���
o ���
o  ����	C  ��          ,���  ����� }��� }���  �����  ��          ,��  ���� ���G ���G  ����  ��          ,��7  ����7 }��c }��c  ����7  ��          ,��� E��� ��� ��� E��� E          ,��'C ���'C ���(o ���(o ���'C �          ,��# E��# ���O ���O E��# E          ,��-� ���-� ���.� ���.� ���-� �          ,��7� E��7� ���8� ���8� E��7� E          ,��#� E��#� ���%' ���%' E��#� E          ,��,� E��,� ���.� ���.� E��,� E          ,��	� ���	� ���
� ���
� ���	� �          ,��:� ���:� ���<� ���<� ���:� �          ,��7� }��7� E��9O E��9O }��7� }          ,��(� }��(� E��0� E��0� }��(� }          ,�� E�� ���/ ���/ E�� E          ,��1 ���1 ���2� ���2� ���1 �          ,��#� }��#� E��&� E��&� }��#� }          ,��� ���� ���� ���� ���� �          ,��k ���k ��� ; ��� ; ���k �          ,��7 }��7 E��� E��� }��7 }          ,�� ��� ���� ���� ��� �          ,��� }��� E��/ E��/ }��� }          ,��	C ���	C ���
� ���
� ���	C �          ,��� ���� ���8� ���8� ���� �          ,���  �����  ����2�  ����2�  �����  ��          ,��'C ���'C ���.� ���.� ���'C �          ,�� E�� ���# ���# E�� E          ,��:� O��:� ���<� ���<� O��:� O          ,��	C O��	C ���
� ���
� O��	C O      !    ,��? ��? ���	 ���	 ��?       !    ,��? +��? ��	 ��	 +��? +      !    ,��? 	7��? 
��	 
��	 	7��? 	7      !    ,��� ��� ���c ���c ���       !    ,��� +��� ��c ��c +��� +      !    ,��� 	7��� 
��c 
��c 	7��� 	7      !    ,��� ��� ���� ���� ���       !    ,��� +��� ��� ��� +��� +      !    ,��� 	7��� 
��� 
��� 	7��� 	7      !    ,��6/ ��6/ ���7 ���7 ��6/       !    ,��6/ +��6/ ��7 ��7 +��6/ +      !    ,��6/ 	7��6/ 
��7 
��7 	7��6/ 	7      !    ,��9w ��9w ���:S ���:S ��9w       !    ,��9w +��9w ��:S ��:S +��9w +      !    ,��9w 	7��9w 
��:S 
��:S 	7��9w 	7      !    ,��<� ��<� ���=� ���=� ��<�       !    ,��<� +��<� ��=� ��=� +��<� +      !    ,��<� 	7��<� 
��=� 
��=� 	7��<� 	7      !    ,��" ��" ���#[ ���#[ ��"       !    ,��" +��" ��#[ ��#[ +��" +      !    ,��" 	7��" 
��#[ 
��#[ 	7��" 	7      !    ,��%� ��%� ���&� ���&� ��%�       !    ,��%� +��%� ��&� ��&� +��%� +      !    ,��%� 	7��%� 
��&� 
��&� 	7��%� 	7      !    ,��) ��) ���)� ���)� ��)       !    ,��) +��) ��)� ��)� +��) +      !    ,��) 	7��) 
��)� 
��)� 	7��) 	7      !    ,��,W ��,W ���-3 ���-3 ��,W       !    ,��,W +��,W ��-3 ��-3 +��,W +      !    ,��,W 	7��,W 
��-3 
��-3 	7��,W 	7      !    ,��/� ��/� ���0{ ���0{ ��/�       !    ,��/� +��/� ��0{ ��0{ +��/� +      !    ,��/� 	7��/� 
��0{ 
��0{ 	7��/� 	7      !    ,��2� ��2� ���3� ���3� ��2�       !    ,��2� +��2� ��3� ��3� +��2� +      !    ,��2� 	7��2� 
��3� 
��3� 	7��2� 	7      !    ,��� 	7��� 
��� 
��� 	7��� 	7      !    ,��� +��� ��� ��� +��� +      !    ,��� ��� ���� ���� ���       !    ,��� 	7��� 
��� 
��� 	7��� 	7      !    ,��� +��� ��� ��� +��� +      !    ,��� ��� ���� ���� ���       !    ,��_ 	7��_ 
��; 
��; 	7��_ 	7      !    ,��_ +��_ ��; ��; +��_ +      !    ,��_ ��_ ���; ���; ��_       !    ,�� 	7�� 
��� 
��� 	7�� 	7      !    ,�� +�� ��� ��� +�� +      !    ,�� �� ���� ���� ��       !    ,��7 	7��7 
��  
��  	7��7 	7      !    ,��7 +��7 ��  ��  +��7 +      !    ,��7 ��7 ���  ���  ��7       !    ,��� ���� ���� ���� ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��W ���W ���3 ���3 ���W �      !    ,��� ���� ���{ ���{ ���� �      !    ,�� ��� ���� ���� ��� �      !    ,��K ���K ���' ���' ���K �      !    ,��� ���� ���o ���o ���� �      !    ,�� � ��� � ���!� ���!� ��� � �      !    ,��$# ���$# ���$� ���$� ���$# �      !    ,��'k ���'k ���(G ���(G ���'k �      !    ,��*� ���*� ���+� ���+� ���*� �      !    ,��6� ���6� ���7� ���7� ���6� �      !    ,��9� ���9� ���:� ���:� ���9� �      !    ,��=7 ���=7 ���> ���> ���=7 �      !    ,��-� ���-� ���.� ���.� ���-� �      !    ,��3_ ���3_ ���4; ���4; ���3_ �      !    ,��" ���" x��#[ x��#[ ���" �      !    ,��� ���� x��� x��� ���� �      !    ,�� ��� x��� x��� ��� �      !    ,��o ���o x��K x��K ���o �      !    ,��� ���� x��� x��� ���� �      !    ,�� ��� x��� x��� ��� �      !    ,��9� ���9� x��:� x��:� ���9� �      !    ,��5? ���5? x��6 x��6 ���5? �      !    ,��0� ���0� x��1k x��1k ���0� �      !    ,��+� ���+� x��,� x��,� ���+� �      !    ,��'/ ���'/ x��( x��( ���'/ �      !    ,��"  ���"  ����#[  ����#[  ���"  �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,��o  ���o  ����K  ����K  ���o  �      !    ,���  ����  �����  �����  ����  �      !    ,��  ���  �����  �����  ���  �      !    ,��9�  ���9�  ����:�  ����:�  ���9�  �      !    ,��5?  ���5?  ����6  ����6  ���5?  �      !    ,��0�  ���0�  ����1k  ����1k  ���0�  �      !    ,��+�  ���+�  ����,�  ����,�  ���+�  �      !    ,��'/  ���'/  ����(  ����(  ���'/  �      !    ,��;W ���;W ���<3 ���<3 ���;W �      !    ,��-. ���-. ���.
 ���.
 ���-. �      !    ,��	� ���	� ���
� ���
� ���	� �      !    ,��� ���� ���� ���� ���� �   	   "    !     4��=� &��=� o��>1 o��>1 ���=- ���=- i   	   "    !     $��8 x��8 k��� k��� !   	   "    !     4��5 ��5 o��� o��� ���� ���� i   	   "    !     $��6� x��6� k��7 k��7 !   	   "    !     $��.i !��.i o��0 o��0 i   	   "    !     $��q !��q o��� o��� i   	   "    !     ��"� 	Z��"� i   	   "    !    � ��; ���
� �   	   "    !    � ��;  ����
�  ��   	   "    !     ��} o��}  �!   	   "    !     �� o��  �!   	   "    !     ��'� o��'�  �!   	   "    !     ��3� o��3�  �!   	   "    !     ��:] o��:]  �!   	   "    !     ��� ���� i   	   "    !     ��� ���� i   	   "    !     �� ��� i   	   "    !     ��,� ���,� i   	   "    !     ��3U ���3U i   	   "    !     ��9� ���9� i   	   "    !     $��] ���] f��&5 f��&5 i   	   "    !     $��� o���  ����$�  ����$� o   	   "    !     $��!I ���!I c��+! c��+! !      "    ,��(o ���(o ���*� ���*� ���(o �      "    ,��� ���� ��� � ��� � ���� �      "    ,��� ?��� y�� y�� ?��� ?      "    ,��-[  ���-[ ���0� ���0�  ���-[  �      "    ,��:� O��:� H��<� H��<� O��:� O      "    ,��6 E��6 ���7� ���7� E��6 E      "    ,��,� E��,� ���.� ���.� E��,� E      "    ,��=� ���=� ���?� ���?� ���=� �      "    ,��( ���( ��� ��� ���( �      "    ,��	C O��	C /��
� /��
� O��	C O      "    ,��7  ���7 ��� ���  ���7  �      "    ,��> }��> ���� ���� }��> }      "    ,��� E��� ���� ���� E��� E          ,��� ���� m��?� m��?� ���� �      #    ,��# 	#��# 
'�� ' 
'�� ' 	#��# 	#      #    ,��# ��# �� ' �� ' ��#       #    ,��# ��# �� ' �� ' ��#       #    ,��(� ��(� ��)� ��)� ��(�       #    ,��(� ��(� ��)� ��)� ��(�       #    ,��(� 	#��(� 
'��)� 
'��)� 	#��(� 	#      #    ,�� ��� ���� ���� ��� �      #    ,��/1 ���/1 ���05 ���05 ���/1 �      #    ,��;C ���;C ���<G ���<G ���;C �      #    ,��6\ ��6\ ��7` ��7` ��6\       #    ,��- ���- ���. ���. ���- �      #    ,��>; ���>; ���?? ���?? ���>; �      #    ,��� ���� ���� ���� ���� �      #    ,��	� ���	� ���
� ���
� ���	� �      #    ,��� ���� ���� ���� ���� �      #    ,��u ��u ��y ��y ��u       #    ,��� ���� ���� ���� ���� �   	   $    !    , ��.} 5��< 5��< %   	   $    !    , ��-8 ���7 �   	   $    !    , ��� 5��	� 5��	� %   	   $    !    , �� ���    	   $    !    , ��- ���)� �   	   $    !    , �� v�� U      $    ,��(o ���(o ���*� ���*� ���(o �      $    ,��� ���� ��� � ��� � ���� �      $    ,��� ?��� y�� y�� ?��� ?      $    ,��-[  ���-[ ���0� ���0�  ���-[  �      $    ,��6 E��6 ���7� ���7� E��6 E      $    ,��,� E��,� ���.� ���.� E��,� E      $    ,��=� ���=� ���?� ���?� ���=� �      $    ,��( ���( ��� ��� ���( �      $    ,��	C O��	C /��
� /��
� O��	C O      $    ,��7  ���7 ��� ���  ���7  �      $    ,��> }��> ���� ���� }��> }      $    ,��� E��� ���O ���O E��� E      $    ,��:� O��:� H��<� H��<� O��:� O          ,��� G��� ���>; ���>; G��� G          ,��	�  ����	�  �a��<$  �a��<$  ����	�  ��           ,��	� )��	� ���<$ ���<$ )��	� )           ,��'  ���' ���>� ���>�  ���'  �      $  
   ��� � L       $  
   ��� J E       $  
   ��? x G       "  
   ��7�  VDD       "  
   ��7�  �� VSS       