magic
tech gf180mcuD
timestamp 1755595969
<< nwell >>
rect 0 63 392 127
rect 0 -99 392 -49
rect 18 -113 373 -99
<< nmos >>
rect 19 21 25 38
rect 36 21 42 38
rect 49 21 55 38
rect 72 21 78 38
rect 85 21 91 38
rect 102 21 108 38
rect 149 21 155 38
rect 166 21 172 38
rect 199 21 205 38
rect 216 21 222 38
rect 227 21 233 38
rect 244 21 250 38
rect 277 21 283 38
rect 294 21 300 38
rect 310 21 316 38
rect 333 21 339 38
rect 349 21 355 38
rect 366 21 372 38
rect 37 -24 43 -7
rect 54 -24 60 -7
rect 70 -24 76 -7
rect 93 -24 99 -7
rect 109 -24 115 -7
rect 126 -24 132 -7
rect 159 -24 165 -7
rect 176 -24 182 -7
rect 187 -24 193 -7
rect 204 -24 210 -7
rect 237 -24 243 -7
rect 254 -24 260 -7
rect 316 -24 322 -7
rect 333 -24 339 -7
<< pmos >>
rect 19 72 25 106
rect 36 72 42 106
rect 49 72 55 106
rect 72 72 78 106
rect 85 72 91 106
rect 102 72 108 106
rect 135 72 141 106
rect 152 72 158 106
rect 163 72 169 106
rect 180 72 186 106
rect 213 72 219 106
rect 230 72 236 106
rect 277 72 283 106
rect 294 72 300 106
rect 310 72 316 106
rect 333 72 339 106
rect 349 72 355 106
rect 366 72 372 106
rect 37 -92 43 -58
rect 54 -92 60 -58
rect 70 -92 76 -58
rect 93 -92 99 -58
rect 109 -92 115 -58
rect 126 -92 132 -58
rect 173 -92 179 -58
rect 190 -92 196 -58
rect 223 -92 229 -58
rect 240 -92 246 -58
rect 251 -92 257 -58
rect 268 -92 274 -58
rect 302 -92 308 -58
rect 319 -92 325 -58
rect 330 -92 336 -58
rect 347 -92 353 -58
<< ndiff >>
rect 58 38 68 39
rect 9 36 19 38
rect 9 23 11 36
rect 16 23 19 36
rect 9 21 19 23
rect 25 36 36 38
rect 25 23 28 36
rect 33 23 36 36
rect 25 21 36 23
rect 42 21 49 38
rect 55 37 72 38
rect 55 23 61 37
rect 66 23 72 37
rect 55 21 72 23
rect 78 21 85 38
rect 91 36 102 38
rect 91 23 94 36
rect 99 23 102 36
rect 91 21 102 23
rect 108 36 118 38
rect 108 23 111 36
rect 116 23 118 36
rect 108 21 118 23
rect 139 36 149 38
rect 139 23 141 36
rect 146 23 149 36
rect 139 21 149 23
rect 155 36 166 38
rect 155 23 158 36
rect 163 23 166 36
rect 155 21 166 23
rect 172 36 182 38
rect 172 23 175 36
rect 180 23 182 36
rect 172 21 182 23
rect 188 32 199 38
rect 188 26 190 32
rect 196 26 199 32
rect 188 21 199 26
rect 205 29 216 38
rect 205 23 208 29
rect 213 23 216 29
rect 205 21 216 23
rect 222 21 227 38
rect 233 36 244 38
rect 233 23 236 36
rect 241 23 244 36
rect 233 21 244 23
rect 250 32 261 38
rect 250 26 253 32
rect 259 26 261 32
rect 250 21 261 26
rect 267 36 277 38
rect 267 23 269 36
rect 274 23 277 36
rect 267 21 277 23
rect 283 36 294 38
rect 283 23 286 36
rect 291 23 294 36
rect 283 21 294 23
rect 300 21 310 38
rect 316 28 333 38
rect 316 23 322 28
rect 327 23 333 28
rect 316 21 333 23
rect 339 21 349 38
rect 355 35 366 38
rect 355 23 358 35
rect 363 23 366 35
rect 355 21 366 23
rect 372 36 382 38
rect 372 23 375 36
rect 380 23 382 36
rect 372 21 382 23
rect 27 -9 37 -7
rect 27 -22 29 -9
rect 34 -22 37 -9
rect 27 -24 37 -22
rect 43 -9 54 -7
rect 43 -22 46 -9
rect 51 -22 54 -9
rect 43 -24 54 -22
rect 60 -24 70 -7
rect 76 -9 93 -7
rect 76 -14 82 -9
rect 87 -14 93 -9
rect 76 -24 93 -14
rect 99 -24 109 -7
rect 115 -9 126 -7
rect 115 -21 118 -9
rect 123 -21 126 -9
rect 115 -24 126 -21
rect 132 -9 142 -7
rect 132 -22 135 -9
rect 140 -22 142 -9
rect 132 -24 142 -22
rect 148 -12 159 -7
rect 148 -18 150 -12
rect 156 -18 159 -12
rect 148 -24 159 -18
rect 165 -9 176 -7
rect 165 -15 168 -9
rect 173 -15 176 -9
rect 165 -24 176 -15
rect 182 -24 187 -7
rect 193 -9 204 -7
rect 193 -22 196 -9
rect 201 -22 204 -9
rect 193 -24 204 -22
rect 210 -12 221 -7
rect 210 -18 213 -12
rect 219 -18 221 -12
rect 210 -24 221 -18
rect 227 -9 237 -7
rect 227 -22 229 -9
rect 234 -22 237 -9
rect 227 -24 237 -22
rect 243 -9 254 -7
rect 243 -22 246 -9
rect 251 -22 254 -9
rect 243 -24 254 -22
rect 260 -9 270 -7
rect 260 -22 263 -9
rect 268 -22 270 -9
rect 260 -24 270 -22
rect 306 -9 316 -7
rect 306 -22 308 -9
rect 313 -22 316 -9
rect 306 -24 316 -22
rect 322 -9 333 -7
rect 322 -22 325 -9
rect 330 -22 333 -9
rect 322 -24 333 -22
rect 339 -9 349 -7
rect 339 -22 342 -9
rect 347 -22 349 -9
rect 339 -24 349 -22
<< pdiff >>
rect 9 104 19 106
rect 9 96 11 104
rect 16 96 19 104
rect 9 72 19 96
rect 25 104 36 106
rect 25 96 28 104
rect 33 96 36 104
rect 25 72 36 96
rect 42 72 49 106
rect 55 104 72 106
rect 55 96 61 104
rect 66 96 72 104
rect 55 72 72 96
rect 78 72 85 106
rect 91 104 102 106
rect 91 96 94 104
rect 99 96 102 104
rect 91 72 102 96
rect 108 104 118 106
rect 108 96 111 104
rect 116 96 118 104
rect 108 72 118 96
rect 124 103 135 106
rect 124 97 126 103
rect 132 97 135 103
rect 124 72 135 97
rect 141 104 152 106
rect 141 74 144 104
rect 149 74 152 104
rect 141 72 152 74
rect 158 72 163 106
rect 169 104 180 106
rect 169 81 172 104
rect 177 81 180 104
rect 169 72 180 81
rect 186 103 197 106
rect 186 97 189 103
rect 195 97 197 103
rect 186 72 197 97
rect 203 104 213 106
rect 203 74 205 104
rect 210 74 213 104
rect 203 72 213 74
rect 219 104 230 106
rect 219 79 222 104
rect 227 79 230 104
rect 219 72 230 79
rect 236 104 246 106
rect 236 74 239 104
rect 244 74 246 104
rect 236 72 246 74
rect 267 104 277 106
rect 267 74 269 104
rect 274 74 277 104
rect 267 72 277 74
rect 283 104 294 106
rect 283 80 286 104
rect 291 80 294 104
rect 283 72 294 80
rect 300 72 310 106
rect 316 104 333 106
rect 316 99 322 104
rect 327 99 333 104
rect 316 72 333 99
rect 339 72 349 106
rect 355 104 366 106
rect 355 80 358 104
rect 363 80 366 104
rect 355 72 366 80
rect 372 104 382 106
rect 372 74 375 104
rect 380 74 382 104
rect 372 72 382 74
rect 27 -60 37 -58
rect 27 -90 29 -60
rect 34 -90 37 -60
rect 27 -92 37 -90
rect 43 -66 54 -58
rect 43 -90 46 -66
rect 51 -90 54 -66
rect 43 -92 54 -90
rect 60 -92 70 -58
rect 76 -85 93 -58
rect 76 -90 82 -85
rect 87 -90 93 -85
rect 76 -92 93 -90
rect 99 -92 109 -58
rect 115 -66 126 -58
rect 115 -90 118 -66
rect 123 -90 126 -66
rect 115 -92 126 -90
rect 132 -60 142 -58
rect 132 -90 135 -60
rect 140 -90 142 -60
rect 132 -92 142 -90
rect 163 -60 173 -58
rect 163 -90 165 -60
rect 170 -90 173 -60
rect 163 -92 173 -90
rect 179 -65 190 -58
rect 179 -90 182 -65
rect 187 -90 190 -65
rect 179 -92 190 -90
rect 196 -60 206 -58
rect 196 -90 199 -60
rect 204 -90 206 -60
rect 196 -92 206 -90
rect 212 -83 223 -58
rect 212 -89 214 -83
rect 220 -89 223 -83
rect 212 -92 223 -89
rect 229 -60 240 -58
rect 229 -90 232 -60
rect 237 -90 240 -60
rect 229 -92 240 -90
rect 246 -92 251 -58
rect 257 -67 268 -58
rect 257 -90 260 -67
rect 265 -90 268 -67
rect 257 -92 268 -90
rect 274 -83 285 -58
rect 274 -89 277 -83
rect 283 -89 285 -83
rect 274 -92 285 -89
rect 291 -83 302 -58
rect 291 -89 293 -83
rect 299 -89 302 -83
rect 291 -92 302 -89
rect 308 -60 319 -58
rect 308 -90 311 -60
rect 316 -90 319 -60
rect 308 -92 319 -90
rect 325 -92 330 -58
rect 336 -67 347 -58
rect 336 -90 339 -67
rect 344 -90 347 -67
rect 336 -92 347 -90
rect 353 -83 364 -58
rect 353 -89 356 -83
rect 362 -89 364 -83
rect 353 -92 364 -89
<< ndiffc >>
rect 11 23 16 36
rect 28 23 33 36
rect 61 23 66 37
rect 94 23 99 36
rect 111 23 116 36
rect 141 23 146 36
rect 158 23 163 36
rect 175 23 180 36
rect 190 26 196 32
rect 208 23 213 29
rect 236 23 241 36
rect 253 26 259 32
rect 269 23 274 36
rect 286 23 291 36
rect 322 23 327 28
rect 358 23 363 35
rect 375 23 380 36
rect 29 -22 34 -9
rect 46 -22 51 -9
rect 82 -14 87 -9
rect 118 -21 123 -9
rect 135 -22 140 -9
rect 150 -18 156 -12
rect 168 -15 173 -9
rect 196 -22 201 -9
rect 213 -18 219 -12
rect 229 -22 234 -9
rect 246 -22 251 -9
rect 263 -22 268 -9
rect 308 -22 313 -9
rect 325 -22 330 -9
rect 342 -22 347 -9
<< pdiffc >>
rect 11 96 16 104
rect 28 96 33 104
rect 61 96 66 104
rect 94 96 99 104
rect 111 96 116 104
rect 126 97 132 103
rect 144 74 149 104
rect 172 81 177 104
rect 189 97 195 103
rect 205 74 210 104
rect 222 79 227 104
rect 239 74 244 104
rect 269 74 274 104
rect 286 80 291 104
rect 322 99 327 104
rect 358 80 363 104
rect 375 74 380 104
rect 29 -90 34 -60
rect 46 -90 51 -66
rect 82 -90 87 -85
rect 118 -90 123 -66
rect 135 -90 140 -60
rect 165 -90 170 -60
rect 182 -90 187 -65
rect 199 -90 204 -60
rect 214 -89 220 -83
rect 232 -90 237 -60
rect 260 -90 265 -67
rect 277 -89 283 -83
rect 293 -89 299 -83
rect 311 -90 316 -60
rect 339 -90 344 -67
rect 356 -89 362 -83
<< psubdiff >>
rect 23 10 38 12
rect 23 4 28 10
rect 33 4 38 10
rect 23 2 38 4
rect 57 10 72 12
rect 57 4 62 10
rect 67 4 72 10
rect 57 2 72 4
rect 89 10 104 12
rect 89 4 94 10
rect 99 4 104 10
rect 89 2 104 4
rect 113 10 128 12
rect 113 4 118 10
rect 123 4 128 10
rect 113 2 128 4
rect 136 10 151 12
rect 136 4 141 10
rect 146 4 151 10
rect 136 2 151 4
rect 170 10 185 12
rect 170 4 175 10
rect 180 4 185 10
rect 170 2 185 4
rect 191 10 206 12
rect 191 4 196 10
rect 201 4 206 10
rect 191 2 206 4
rect 228 10 243 12
rect 228 4 233 10
rect 238 4 243 10
rect 228 2 243 4
rect 258 10 273 12
rect 258 4 263 10
rect 268 4 273 10
rect 258 2 273 4
rect 303 10 318 12
rect 303 4 308 10
rect 313 4 318 10
rect 303 2 318 4
rect 337 10 352 12
rect 337 4 342 10
rect 347 4 352 10
rect 337 2 352 4
rect 367 10 382 12
rect 367 4 372 10
rect 377 4 382 10
rect 367 2 382 4
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
rect 54 120 69 122
rect 54 115 59 120
rect 64 115 69 120
rect 54 113 69 115
rect 78 120 93 122
rect 78 115 83 120
rect 88 115 93 120
rect 78 113 93 115
rect 102 120 117 122
rect 102 115 107 120
rect 112 115 117 120
rect 102 113 117 115
rect 136 120 151 122
rect 136 115 141 120
rect 146 115 151 120
rect 136 113 151 115
rect 160 120 175 122
rect 160 115 165 120
rect 170 115 175 120
rect 160 113 175 115
rect 200 120 215 122
rect 200 115 205 120
rect 210 115 215 120
rect 200 113 215 115
rect 224 120 239 122
rect 224 115 229 120
rect 234 115 239 120
rect 224 113 239 115
rect 264 120 279 122
rect 264 115 269 120
rect 274 115 279 120
rect 264 113 279 115
rect 288 120 303 122
rect 288 115 293 120
rect 298 115 303 120
rect 288 113 303 115
rect 312 120 327 122
rect 312 115 317 120
rect 322 115 327 120
rect 312 113 327 115
rect 336 120 351 122
rect 336 115 341 120
rect 346 115 351 120
rect 336 113 351 115
rect 360 120 375 122
rect 360 115 365 120
rect 370 115 375 120
rect 360 113 375 115
rect 24 -101 39 -99
rect 24 -106 29 -101
rect 34 -106 39 -101
rect 24 -108 39 -106
rect 48 -101 63 -99
rect 48 -106 53 -101
rect 58 -106 63 -101
rect 48 -108 63 -106
rect 72 -101 87 -99
rect 72 -106 77 -101
rect 82 -106 87 -101
rect 72 -108 87 -106
rect 96 -101 111 -99
rect 96 -106 101 -101
rect 106 -106 111 -101
rect 96 -108 111 -106
rect 120 -101 135 -99
rect 120 -106 125 -101
rect 130 -106 135 -101
rect 120 -108 135 -106
rect 160 -101 175 -99
rect 160 -106 165 -101
rect 170 -106 175 -101
rect 160 -108 175 -106
rect 184 -101 199 -99
rect 184 -106 189 -101
rect 194 -106 199 -101
rect 184 -108 199 -106
rect 224 -101 239 -99
rect 224 -106 229 -101
rect 234 -106 239 -101
rect 224 -108 239 -106
rect 248 -101 263 -99
rect 248 -106 253 -101
rect 258 -106 263 -101
rect 248 -108 263 -106
rect 303 -101 318 -99
rect 303 -106 308 -101
rect 313 -106 318 -101
rect 303 -108 318 -106
rect 327 -101 342 -99
rect 327 -106 332 -101
rect 337 -106 342 -101
rect 327 -108 342 -106
<< psubdiffcont >>
rect 28 4 33 10
rect 62 4 67 10
rect 94 4 99 10
rect 118 4 123 10
rect 141 4 146 10
rect 175 4 180 10
rect 196 4 201 10
rect 233 4 238 10
rect 263 4 268 10
rect 308 4 313 10
rect 342 4 347 10
rect 372 4 377 10
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
rect 59 115 64 120
rect 83 115 88 120
rect 107 115 112 120
rect 141 115 146 120
rect 165 115 170 120
rect 205 115 210 120
rect 229 115 234 120
rect 269 115 274 120
rect 293 115 298 120
rect 317 115 322 120
rect 341 115 346 120
rect 365 115 370 120
rect 29 -106 34 -101
rect 53 -106 58 -101
rect 77 -106 82 -101
rect 101 -106 106 -101
rect 125 -106 130 -101
rect 165 -106 170 -101
rect 189 -106 194 -101
rect 229 -106 234 -101
rect 253 -106 258 -101
rect 308 -106 313 -101
rect 332 -106 337 -101
<< polysilicon >>
rect 19 106 25 111
rect 36 106 42 111
rect 49 106 55 111
rect 72 106 78 111
rect 85 106 91 111
rect 102 106 108 111
rect 135 106 141 111
rect 152 106 158 111
rect 163 106 169 111
rect 180 106 186 111
rect 213 106 219 111
rect 230 106 236 111
rect 277 106 283 111
rect 294 106 300 111
rect 310 106 316 111
rect 333 106 339 111
rect 349 106 355 111
rect 366 106 372 111
rect 19 54 25 72
rect 36 70 42 72
rect 31 68 42 70
rect 31 62 33 68
rect 39 62 42 68
rect 31 60 42 62
rect 49 70 55 72
rect 72 70 78 72
rect 85 70 91 72
rect 102 70 108 72
rect 49 68 63 70
rect 49 62 55 68
rect 61 62 63 68
rect 49 60 63 62
rect 70 68 80 70
rect 70 62 72 68
rect 78 62 80 68
rect 85 65 108 70
rect 70 60 80 62
rect 19 52 35 54
rect 19 46 27 52
rect 33 51 35 52
rect 33 46 42 51
rect 19 44 42 46
rect 19 38 25 44
rect 36 38 42 44
rect 49 38 55 60
rect 102 54 108 65
rect 135 68 141 72
rect 152 68 158 72
rect 135 63 158 68
rect 163 69 169 72
rect 163 67 172 69
rect 180 67 186 72
rect 163 65 186 67
rect 163 63 172 65
rect 149 54 155 63
rect 60 52 70 54
rect 91 52 108 54
rect 60 46 62 52
rect 68 46 78 52
rect 91 49 93 52
rect 60 44 78 46
rect 72 38 78 44
rect 85 46 93 49
rect 99 46 108 52
rect 85 44 108 46
rect 141 52 155 54
rect 141 46 144 52
rect 150 46 155 52
rect 141 44 155 46
rect 85 38 91 44
rect 102 38 108 44
rect 149 38 155 44
rect 166 59 172 63
rect 178 61 186 65
rect 178 59 180 61
rect 166 57 180 59
rect 166 38 172 57
rect 213 54 219 72
rect 204 52 219 54
rect 204 46 208 52
rect 214 46 219 52
rect 204 44 219 46
rect 199 40 208 44
rect 213 43 219 44
rect 230 67 236 72
rect 277 70 283 72
rect 294 70 300 72
rect 230 65 244 67
rect 230 59 236 65
rect 242 59 244 65
rect 230 57 244 59
rect 277 65 300 70
rect 310 70 316 72
rect 333 70 339 72
rect 310 68 320 70
rect 230 45 236 57
rect 277 54 283 65
rect 310 63 312 68
rect 318 63 320 68
rect 310 61 320 63
rect 329 68 339 70
rect 329 62 331 68
rect 337 62 339 68
rect 349 70 355 72
rect 366 70 372 72
rect 349 65 372 70
rect 329 60 339 62
rect 277 52 290 54
rect 277 46 282 52
rect 288 46 290 52
rect 230 43 250 45
rect 213 40 222 43
rect 199 38 205 40
rect 216 38 222 40
rect 227 40 250 43
rect 227 38 233 40
rect 244 38 250 40
rect 277 44 290 46
rect 305 48 316 50
rect 277 40 300 44
rect 305 42 307 48
rect 313 42 316 48
rect 305 40 316 42
rect 277 38 283 40
rect 294 38 300 40
rect 310 38 316 40
rect 333 38 339 60
rect 345 58 355 60
rect 345 53 347 58
rect 353 53 355 58
rect 366 54 372 65
rect 345 51 355 53
rect 349 38 355 51
rect 360 52 372 54
rect 360 46 362 52
rect 368 46 372 52
rect 360 44 372 46
rect 366 38 372 44
rect 19 16 25 21
rect 36 16 42 21
rect 49 16 55 21
rect 72 16 78 21
rect 85 16 91 21
rect 102 16 108 21
rect 149 16 155 21
rect 166 16 172 21
rect 199 16 205 21
rect 216 16 222 21
rect 227 16 233 21
rect 244 16 250 21
rect 277 16 283 21
rect 294 16 300 21
rect 310 16 316 21
rect 333 16 339 21
rect 349 16 355 21
rect 366 16 372 21
rect 37 -7 43 -2
rect 54 -7 60 -2
rect 70 -7 76 -2
rect 93 -7 99 -2
rect 109 -7 115 -2
rect 126 -7 132 -2
rect 159 -7 165 -2
rect 176 -7 182 -2
rect 187 -7 193 -2
rect 204 -7 210 -2
rect 237 -7 243 -2
rect 254 -7 260 -2
rect 316 -7 322 -2
rect 333 -7 339 -2
rect 37 -26 43 -24
rect 54 -26 60 -24
rect 70 -26 76 -24
rect 37 -30 60 -26
rect 65 -28 76 -26
rect 37 -32 50 -30
rect 37 -38 42 -32
rect 48 -38 50 -32
rect 65 -34 67 -28
rect 73 -34 76 -28
rect 65 -36 76 -34
rect 37 -40 50 -38
rect 37 -51 43 -40
rect 93 -46 99 -24
rect 109 -37 115 -24
rect 126 -30 132 -24
rect 159 -26 165 -24
rect 176 -26 182 -24
rect 159 -30 168 -26
rect 173 -29 182 -26
rect 187 -26 193 -24
rect 204 -26 210 -24
rect 187 -29 210 -26
rect 173 -30 179 -29
rect 105 -39 115 -37
rect 105 -44 107 -39
rect 113 -44 115 -39
rect 120 -32 132 -30
rect 120 -38 122 -32
rect 128 -38 132 -32
rect 120 -40 132 -38
rect 164 -32 179 -30
rect 164 -38 168 -32
rect 174 -38 179 -32
rect 164 -40 179 -38
rect 105 -46 115 -44
rect 70 -49 80 -47
rect 37 -56 60 -51
rect 37 -58 43 -56
rect 54 -58 60 -56
rect 70 -54 72 -49
rect 78 -54 80 -49
rect 70 -56 80 -54
rect 89 -48 99 -46
rect 89 -54 91 -48
rect 97 -54 99 -48
rect 126 -51 132 -40
rect 89 -56 99 -54
rect 70 -58 76 -56
rect 93 -58 99 -56
rect 109 -56 132 -51
rect 109 -58 115 -56
rect 126 -58 132 -56
rect 173 -58 179 -40
rect 190 -31 210 -29
rect 237 -30 243 -24
rect 190 -43 196 -31
rect 229 -32 243 -30
rect 229 -38 232 -32
rect 238 -38 243 -32
rect 229 -40 243 -38
rect 190 -45 204 -43
rect 190 -51 196 -45
rect 202 -51 204 -45
rect 237 -49 243 -40
rect 254 -43 260 -24
rect 316 -30 322 -24
rect 308 -32 322 -30
rect 308 -38 311 -32
rect 317 -38 322 -32
rect 308 -40 322 -38
rect 254 -45 268 -43
rect 254 -49 260 -45
rect 190 -53 204 -51
rect 190 -58 196 -53
rect 223 -54 246 -49
rect 223 -58 229 -54
rect 240 -58 246 -54
rect 251 -51 260 -49
rect 266 -47 268 -45
rect 266 -51 274 -47
rect 316 -49 322 -40
rect 333 -43 339 -24
rect 333 -45 347 -43
rect 333 -49 339 -45
rect 251 -53 274 -51
rect 251 -55 260 -53
rect 251 -58 257 -55
rect 268 -58 274 -53
rect 302 -54 325 -49
rect 302 -58 308 -54
rect 319 -58 325 -54
rect 330 -51 339 -49
rect 345 -47 347 -45
rect 345 -51 353 -47
rect 330 -53 353 -51
rect 330 -55 339 -53
rect 330 -58 336 -55
rect 347 -58 353 -53
rect 37 -97 43 -92
rect 54 -97 60 -92
rect 70 -97 76 -92
rect 93 -97 99 -92
rect 109 -97 115 -92
rect 126 -97 132 -92
rect 173 -97 179 -92
rect 190 -97 196 -92
rect 223 -97 229 -92
rect 240 -97 246 -92
rect 251 -97 257 -92
rect 268 -97 274 -92
rect 302 -97 308 -92
rect 319 -97 325 -92
rect 330 -97 336 -92
rect 347 -97 353 -92
<< polycontact >>
rect 33 62 39 68
rect 55 62 61 68
rect 72 62 78 68
rect 27 46 33 52
rect 62 46 68 52
rect 93 46 99 52
rect 144 46 150 52
rect 172 59 178 65
rect 208 46 214 52
rect 236 59 242 65
rect 312 63 318 68
rect 331 62 337 68
rect 282 46 288 52
rect 307 42 313 48
rect 347 53 353 58
rect 362 46 368 52
rect 42 -38 48 -32
rect 67 -34 73 -28
rect 107 -44 113 -39
rect 122 -38 128 -32
rect 168 -38 174 -32
rect 72 -54 78 -49
rect 91 -54 97 -48
rect 232 -38 238 -32
rect 196 -51 202 -45
rect 311 -38 317 -32
rect 260 -51 266 -45
rect 339 -51 345 -45
<< metal1 >>
rect 0 120 392 127
rect 0 115 11 120
rect 16 115 35 120
rect 40 115 59 120
rect 64 115 83 120
rect 88 115 107 120
rect 112 115 141 120
rect 146 115 165 120
rect 170 115 205 120
rect 210 115 229 120
rect 234 115 269 120
rect 274 115 293 120
rect 298 115 317 120
rect 322 115 341 120
rect 346 115 365 120
rect 370 115 392 120
rect 0 113 392 115
rect 11 104 16 106
rect 11 68 16 96
rect 28 104 33 113
rect 61 104 66 106
rect 28 94 33 96
rect 60 96 61 97
rect 60 91 66 96
rect 94 104 99 113
rect 94 94 99 96
rect 111 104 116 106
rect 60 83 66 85
rect 111 78 116 96
rect 125 103 133 105
rect 125 97 126 103
rect 132 97 133 103
rect 125 95 133 97
rect 144 104 149 113
rect 124 88 132 90
rect 124 82 125 88
rect 131 82 132 88
rect 124 80 132 82
rect 55 73 116 78
rect 55 68 61 73
rect 11 62 33 68
rect 39 62 48 68
rect 11 36 16 62
rect 42 52 48 62
rect 70 62 72 68
rect 78 62 80 68
rect 55 60 61 62
rect 25 46 27 52
rect 33 46 35 52
rect 42 46 62 52
rect 68 46 70 52
rect 91 46 93 52
rect 99 46 101 52
rect 60 39 66 41
rect 11 21 16 23
rect 28 36 33 38
rect 60 30 61 33
rect 28 14 33 23
rect 61 21 66 23
rect 94 36 99 38
rect 94 14 99 23
rect 111 36 116 73
rect 125 52 131 80
rect 172 104 177 106
rect 188 103 196 105
rect 188 97 189 103
rect 195 97 196 103
rect 188 95 196 97
rect 205 104 210 113
rect 172 79 177 81
rect 158 78 177 79
rect 144 72 149 74
rect 156 72 158 78
rect 164 74 177 78
rect 222 104 227 106
rect 222 78 227 79
rect 239 104 244 113
rect 164 72 166 74
rect 205 72 210 74
rect 220 72 222 78
rect 228 72 230 78
rect 239 72 244 74
rect 269 104 274 106
rect 286 104 291 113
rect 322 104 327 106
rect 322 93 327 99
rect 321 91 327 93
rect 358 104 363 113
rect 319 85 321 91
rect 327 85 329 91
rect 286 78 291 80
rect 125 46 144 52
rect 150 46 152 52
rect 111 21 116 23
rect 141 36 146 38
rect 141 14 146 23
rect 158 36 163 72
rect 170 59 172 65
rect 178 59 180 65
rect 206 46 208 52
rect 214 46 216 52
rect 158 21 163 23
rect 175 36 180 38
rect 222 37 227 72
rect 269 67 274 74
rect 312 75 352 80
rect 358 78 363 80
rect 375 104 380 106
rect 312 68 318 75
rect 347 70 352 75
rect 375 70 380 74
rect 331 68 337 70
rect 234 59 236 65
rect 242 59 244 65
rect 269 62 305 67
rect 310 63 312 68
rect 318 63 320 68
rect 189 32 197 34
rect 189 26 190 32
rect 196 26 197 32
rect 189 24 197 26
rect 208 32 227 37
rect 236 36 241 38
rect 208 29 213 32
rect 175 14 180 23
rect 208 21 213 23
rect 269 36 274 62
rect 299 58 305 62
rect 331 58 337 62
rect 347 64 380 70
rect 347 59 353 64
rect 299 53 337 58
rect 345 58 355 59
rect 345 53 347 58
rect 353 53 355 58
rect 280 46 282 52
rect 288 46 290 52
rect 360 48 362 52
rect 305 42 307 48
rect 313 46 362 48
rect 368 46 370 52
rect 313 42 367 46
rect 252 32 260 34
rect 252 26 253 32
rect 259 26 260 32
rect 252 24 260 26
rect 236 14 241 23
rect 269 21 274 23
rect 286 36 291 38
rect 321 36 327 37
rect 319 30 321 36
rect 327 30 329 36
rect 358 35 363 37
rect 321 28 327 30
rect 286 14 291 23
rect 322 21 327 23
rect 358 14 363 23
rect 375 36 380 64
rect 375 21 380 23
rect 0 10 392 14
rect 0 4 28 10
rect 33 4 62 10
rect 67 4 94 10
rect 99 4 118 10
rect 123 4 141 10
rect 146 4 175 10
rect 180 4 196 10
rect 201 4 233 10
rect 238 4 263 10
rect 268 4 308 10
rect 313 4 342 10
rect 347 4 372 10
rect 377 4 392 10
rect 0 0 392 4
rect 29 -9 34 -7
rect 29 -48 34 -22
rect 46 -9 51 0
rect 82 -9 87 -7
rect 81 -16 87 -14
rect 118 -9 123 0
rect 79 -22 81 -16
rect 87 -22 89 -16
rect 46 -24 51 -22
rect 81 -23 87 -22
rect 118 -23 123 -21
rect 135 -9 140 -7
rect 168 -9 173 -7
rect 149 -12 157 -10
rect 149 -18 150 -12
rect 156 -18 157 -12
rect 149 -20 157 -18
rect 168 -18 173 -15
rect 196 -9 201 0
rect 40 -38 42 -32
rect 48 -38 50 -32
rect 65 -34 67 -28
rect 73 -32 127 -28
rect 73 -34 122 -32
rect 120 -38 122 -34
rect 128 -38 130 -32
rect 59 -44 97 -39
rect 59 -48 65 -44
rect 29 -53 65 -48
rect 91 -48 97 -44
rect 105 -44 107 -39
rect 113 -44 115 -39
rect 105 -45 115 -44
rect 29 -60 34 -53
rect 70 -54 72 -49
rect 78 -54 80 -49
rect 72 -61 78 -54
rect 91 -56 97 -54
rect 107 -50 113 -45
rect 135 -50 140 -22
rect 168 -23 187 -18
rect 166 -38 168 -32
rect 174 -38 176 -32
rect 107 -56 140 -50
rect 107 -61 112 -56
rect 29 -92 34 -90
rect 46 -66 51 -64
rect 72 -66 112 -61
rect 135 -60 140 -56
rect 182 -58 187 -23
rect 229 -9 234 0
rect 212 -12 220 -10
rect 212 -18 213 -12
rect 219 -18 220 -12
rect 212 -20 220 -18
rect 196 -24 201 -22
rect 229 -24 234 -22
rect 246 -9 251 -7
rect 230 -38 232 -32
rect 238 -38 240 -32
rect 194 -51 196 -45
rect 202 -51 204 -45
rect 246 -58 251 -22
rect 263 -9 268 0
rect 263 -24 268 -22
rect 308 -9 313 0
rect 308 -24 313 -22
rect 325 -9 330 -7
rect 309 -38 311 -32
rect 317 -38 319 -32
rect 258 -51 260 -45
rect 266 -51 268 -45
rect 325 -58 330 -22
rect 342 -9 347 0
rect 342 -24 347 -22
rect 337 -51 339 -45
rect 345 -51 347 -45
rect 118 -66 123 -64
rect 79 -77 81 -71
rect 87 -77 89 -71
rect 81 -79 87 -77
rect 46 -99 51 -90
rect 82 -85 87 -79
rect 82 -92 87 -90
rect 118 -99 123 -90
rect 135 -92 140 -90
rect 165 -60 170 -58
rect 180 -64 182 -58
rect 188 -64 190 -58
rect 199 -60 204 -58
rect 165 -99 170 -90
rect 182 -65 187 -64
rect 182 -92 187 -90
rect 232 -60 237 -58
rect 199 -99 204 -90
rect 213 -83 221 -81
rect 213 -89 214 -83
rect 220 -89 221 -83
rect 213 -91 221 -89
rect 244 -64 246 -58
rect 252 -60 254 -58
rect 311 -60 316 -58
rect 252 -64 265 -60
rect 246 -65 265 -64
rect 232 -99 237 -90
rect 260 -67 265 -65
rect 260 -92 265 -90
rect 276 -83 284 -81
rect 276 -89 277 -83
rect 283 -89 284 -83
rect 276 -91 284 -89
rect 292 -83 300 -81
rect 292 -89 293 -83
rect 299 -89 300 -83
rect 292 -91 300 -89
rect 323 -64 325 -58
rect 331 -60 333 -58
rect 331 -64 344 -60
rect 325 -65 344 -64
rect 311 -99 316 -90
rect 339 -67 344 -65
rect 339 -92 344 -90
rect 355 -83 363 -81
rect 355 -89 356 -83
rect 362 -89 363 -83
rect 355 -91 363 -89
rect 0 -101 392 -99
rect 0 -106 29 -101
rect 34 -106 53 -101
rect 58 -106 77 -101
rect 82 -106 101 -101
rect 106 -106 125 -101
rect 130 -106 165 -101
rect 170 -106 189 -101
rect 194 -106 229 -101
rect 234 -106 253 -101
rect 258 -106 308 -101
rect 313 -106 332 -101
rect 337 -106 392 -101
rect 0 -113 392 -106
<< via1 >>
rect 60 85 66 91
rect 126 97 132 103
rect 125 82 131 88
rect 72 62 78 68
rect 27 46 33 52
rect 93 46 99 52
rect 60 37 66 39
rect 60 33 61 37
rect 61 33 66 37
rect 189 97 195 103
rect 158 72 164 78
rect 222 72 228 78
rect 321 85 327 91
rect 144 46 150 52
rect 172 59 178 65
rect 208 46 214 52
rect 236 59 242 65
rect 190 26 196 32
rect 282 46 288 52
rect 362 46 368 52
rect 253 26 259 32
rect 321 30 327 36
rect 81 -22 87 -16
rect 150 -18 156 -12
rect 42 -38 48 -32
rect 122 -38 128 -32
rect 168 -38 174 -32
rect 213 -18 219 -12
rect 232 -38 238 -32
rect 196 -51 202 -45
rect 311 -38 317 -32
rect 260 -51 266 -45
rect 339 -51 345 -45
rect 81 -77 87 -71
rect 182 -64 188 -58
rect 214 -89 220 -83
rect 246 -64 252 -58
rect 277 -89 283 -83
rect 293 -89 299 -83
rect 325 -64 331 -58
rect 356 -89 362 -83
<< metal2 >>
rect 124 103 197 104
rect 124 97 126 103
rect 132 97 189 103
rect 195 97 197 103
rect 60 92 66 97
rect 124 96 197 97
rect 208 97 288 103
rect 59 91 67 92
rect 59 85 60 91
rect 66 90 67 91
rect 208 90 214 97
rect 66 88 132 90
rect 66 85 125 88
rect 59 84 125 85
rect 59 83 66 84
rect 27 53 33 54
rect 26 52 34 53
rect 26 46 27 52
rect 33 46 34 52
rect 26 45 34 46
rect 27 26 33 45
rect 59 40 65 83
rect 124 82 125 84
rect 131 82 132 88
rect 124 80 132 82
rect 158 84 214 90
rect 158 79 166 84
rect 156 78 166 79
rect 156 72 158 78
rect 164 72 166 78
rect 156 71 166 72
rect 220 78 230 79
rect 220 72 222 78
rect 228 72 230 78
rect 220 71 230 72
rect 72 69 79 70
rect 71 68 80 69
rect 71 62 72 68
rect 78 65 150 68
rect 170 65 180 66
rect 78 62 172 65
rect 71 61 80 62
rect 72 60 80 61
rect 58 39 68 40
rect 58 33 60 39
rect 66 33 68 39
rect 58 32 68 33
rect 74 26 80 60
rect 144 59 172 62
rect 178 59 180 65
rect 170 58 180 59
rect 234 58 235 66
rect 243 65 244 66
rect 243 59 274 65
rect 243 58 244 59
rect 93 53 99 54
rect 92 52 100 53
rect 142 52 152 53
rect 206 52 216 53
rect 91 46 93 52
rect 99 46 101 52
rect 142 46 144 52
rect 150 46 208 52
rect 214 46 216 52
rect 92 45 100 46
rect 142 45 152 46
rect 206 45 216 46
rect 93 44 99 45
rect 27 20 80 26
rect 188 32 198 33
rect 251 32 261 33
rect 188 26 190 32
rect 196 26 253 32
rect 259 26 261 32
rect 188 25 198 26
rect 251 25 261 26
rect 268 23 274 59
rect 282 53 288 97
rect 321 92 327 93
rect 320 91 328 92
rect 320 85 321 91
rect 327 85 383 91
rect 320 84 328 85
rect 281 52 289 53
rect 280 46 282 52
rect 288 46 290 52
rect 281 45 289 46
rect 321 37 327 84
rect 361 52 369 53
rect 360 46 362 52
rect 368 46 370 52
rect 361 45 369 46
rect 319 36 329 37
rect 319 30 321 36
rect 327 30 329 36
rect 319 29 329 30
rect 362 23 368 45
rect 268 17 368 23
rect 42 -9 142 -3
rect 42 -31 48 -9
rect 79 -16 89 -15
rect 79 -22 81 -16
rect 87 -22 89 -16
rect 79 -23 89 -22
rect 41 -32 49 -31
rect 40 -38 42 -32
rect 48 -38 50 -32
rect 41 -39 49 -38
rect 81 -70 87 -23
rect 136 -26 142 -9
rect 148 -12 158 -11
rect 211 -12 221 -11
rect 148 -18 150 -12
rect 156 -18 213 -12
rect 219 -18 221 -12
rect 148 -19 158 -18
rect 211 -19 221 -18
rect 136 -31 174 -26
rect 121 -32 129 -31
rect 136 -32 176 -31
rect 120 -38 122 -32
rect 128 -38 130 -32
rect 166 -38 168 -32
rect 174 -38 176 -32
rect 121 -39 129 -38
rect 166 -39 176 -38
rect 230 -32 240 -31
rect 268 -32 274 17
rect 230 -38 232 -32
rect 238 -38 274 -32
rect 309 -32 319 -31
rect 376 -32 383 85
rect 309 -38 311 -32
rect 317 -38 383 -32
rect 230 -39 240 -38
rect 309 -39 319 -38
rect 194 -45 204 -44
rect 258 -45 268 -44
rect 337 -45 347 -44
rect 152 -51 196 -45
rect 202 -51 260 -45
rect 266 -51 268 -45
rect 80 -71 88 -70
rect 152 -71 158 -51
rect 194 -52 204 -51
rect 258 -52 268 -51
rect 293 -51 339 -45
rect 345 -51 347 -45
rect 180 -65 181 -57
rect 189 -65 190 -57
rect 244 -58 254 -57
rect 293 -58 299 -51
rect 337 -52 347 -51
rect 244 -64 246 -58
rect 252 -64 299 -58
rect 323 -58 333 -57
rect 323 -64 325 -58
rect 331 -64 333 -58
rect 244 -65 254 -64
rect 323 -65 333 -64
rect 80 -77 81 -71
rect 87 -77 158 -71
rect 80 -78 88 -77
rect 81 -79 87 -78
rect 212 -83 285 -82
rect 212 -89 214 -83
rect 220 -89 277 -83
rect 283 -89 285 -83
rect 212 -90 285 -89
rect 291 -83 364 -82
rect 291 -89 293 -83
rect 299 -89 356 -83
rect 362 -89 364 -83
rect 291 -90 364 -89
<< via2 >>
rect 235 65 243 66
rect 235 59 236 65
rect 236 59 242 65
rect 242 59 243 65
rect 235 58 243 59
rect 181 -58 189 -57
rect 181 -64 182 -58
rect 182 -64 188 -58
rect 188 -64 189 -58
rect 181 -65 189 -64
<< metal3 >>
rect 234 66 244 67
rect 234 65 235 66
rect 182 59 235 65
rect 182 -56 188 59
rect 234 58 235 59
rect 243 58 244 66
rect 234 57 244 58
rect 180 -57 190 -56
rect 180 -65 181 -57
rect 189 -65 190 -57
rect 180 -66 190 -65
<< labels >>
rlabel metal2 30 49 30 49 1 my_nxor_0.A
rlabel metal2 63 87 63 87 1 my_nxor_0.Y
rlabel metal2 96 49 96 49 1 my_nxor_0.B
rlabel via1 161 75 161 75 1 my_nor_0.Y
rlabel metal2 211 49 211 49 1 my_nand_0.A
rlabel via2 239 62 239 62 1 my_nand_0.B
rlabel metal2 225 75 225 75 1 my_nand_0.Y
rlabel via1 84 -73 84 -73 5 my_xor_0.Y
rlabel via1 125 -35 125 -35 5 my_xor_0.B
rlabel via1 45 -35 45 -35 5 my_xor_0.A
rlabel via1 235 -35 235 -35 1 my_nor_1.A
rlabel via1 263 -48 263 -48 1 my_nor_1.B
rlabel via1 249 -61 249 -61 1 my_nor_1.Y
rlabel via1 314 -35 314 -35 1 my_nor_2.A
rlabel via1 342 -48 342 -48 1 my_nor_2.B
rlabel via1 328 -61 328 -61 1 my_nor_2.Y
rlabel via1 285 49 285 49 1 my_xor_1.A
rlabel via1 365 49 365 49 1 my_xor_1.B
rlabel via1 324 88 324 88 1 my_xor_1.Y
rlabel via1 171 -35 171 -35 1 my_nand_1.A
rlabel via1 199 -48 199 -48 1 my_nand_1.B
rlabel via1 185 -61 185 -61 1 my_nand_1.Y
rlabel metal1 3 -106 3 -106 1 VDD
rlabel metal1 4 121 4 121 1 VDD
rlabel metal1 4 7 4 7 1 VSS
rlabel via1 30 47 30 47 1 B1
rlabel via1 96 47 96 47 1 A1
rlabel via1 45 -34 45 -34 1 B0
rlabel via1 125 -34 125 -34 1 A0
rlabel via1 147 49 147 49 1 my_nor_0.B
rlabel via1 175 62 175 62 1 my_nor_0.A
rlabel via1 324 87 324 87 1 L
rlabel via1 328 -63 328 -63 1 G
rlabel via1 249 -63 249 -63 1 E
<< end >>
