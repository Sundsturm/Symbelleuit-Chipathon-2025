magic
tech gf180mcuD
magscale 1 10
timestamp 1757081687
<< nwell >>
rect -12807 13441 -9831 14153
<< nmos >>
rect -12633 13139 -12573 13309
rect -12465 13139 -12405 13309
rect -12129 13139 -12069 13309
rect -12021 13139 -11961 13309
rect -11685 13139 -11625 13309
rect -11517 13139 -11457 13309
rect -11181 13139 -11121 13309
rect -11013 13139 -10953 13309
rect -10677 13139 -10617 13309
rect -10569 13139 -10509 13309
rect -10233 13139 -10173 13309
rect -10065 13139 -10005 13309
<< pmos >>
rect -12609 13531 -12549 13871
rect -12441 13531 -12381 13871
rect -12105 13531 -12045 13871
rect -11937 13531 -11877 13871
rect -11769 13531 -11709 13871
rect -11601 13531 -11541 13871
rect -11265 13531 -11205 13871
rect -11097 13531 -11037 13871
rect -10761 13531 -10701 13871
rect -10593 13531 -10533 13871
rect -10257 13531 -10197 13871
rect -10089 13531 -10029 13871
<< ndiff >>
rect -12741 13247 -12633 13309
rect -12741 13201 -12710 13247
rect -12664 13201 -12633 13247
rect -12741 13139 -12633 13201
rect -12573 13247 -12465 13309
rect -12573 13201 -12542 13247
rect -12496 13201 -12465 13247
rect -12573 13139 -12465 13201
rect -12405 13247 -12297 13309
rect -12405 13201 -12374 13247
rect -12328 13201 -12297 13247
rect -12405 13139 -12297 13201
rect -12237 13247 -12129 13309
rect -12237 13201 -12206 13247
rect -12160 13201 -12129 13247
rect -12237 13139 -12129 13201
rect -12069 13139 -12021 13309
rect -11961 13247 -11853 13309
rect -11961 13201 -11930 13247
rect -11884 13201 -11853 13247
rect -11961 13139 -11853 13201
rect -11793 13247 -11685 13309
rect -11793 13201 -11762 13247
rect -11716 13201 -11685 13247
rect -11793 13139 -11685 13201
rect -11625 13247 -11517 13309
rect -11625 13201 -11594 13247
rect -11548 13201 -11517 13247
rect -11625 13139 -11517 13201
rect -11457 13247 -11349 13309
rect -11457 13201 -11426 13247
rect -11380 13201 -11349 13247
rect -11457 13139 -11349 13201
rect -11289 13247 -11181 13309
rect -11289 13201 -11258 13247
rect -11212 13201 -11181 13247
rect -11289 13139 -11181 13201
rect -11121 13247 -11013 13309
rect -11121 13201 -11090 13247
rect -11044 13201 -11013 13247
rect -11121 13139 -11013 13201
rect -10953 13247 -10845 13309
rect -10953 13201 -10922 13247
rect -10876 13201 -10845 13247
rect -10953 13139 -10845 13201
rect -10785 13247 -10677 13309
rect -10785 13201 -10754 13247
rect -10708 13201 -10677 13247
rect -10785 13139 -10677 13201
rect -10617 13139 -10569 13309
rect -10509 13247 -10401 13309
rect -10509 13201 -10478 13247
rect -10432 13201 -10401 13247
rect -10509 13139 -10401 13201
rect -10341 13247 -10233 13309
rect -10341 13201 -10310 13247
rect -10264 13201 -10233 13247
rect -10341 13139 -10233 13201
rect -10173 13247 -10065 13309
rect -10173 13201 -10142 13247
rect -10096 13201 -10065 13247
rect -10173 13139 -10065 13201
rect -10005 13247 -9897 13309
rect -10005 13201 -9974 13247
rect -9928 13201 -9897 13247
rect -10005 13139 -9897 13201
<< pdiff >>
rect -12717 13818 -12609 13871
rect -12717 13584 -12686 13818
rect -12640 13584 -12609 13818
rect -12717 13531 -12609 13584
rect -12549 13818 -12441 13871
rect -12549 13584 -12518 13818
rect -12472 13584 -12441 13818
rect -12549 13531 -12441 13584
rect -12381 13818 -12273 13871
rect -12381 13584 -12350 13818
rect -12304 13584 -12273 13818
rect -12381 13531 -12273 13584
rect -12213 13818 -12105 13871
rect -12213 13584 -12182 13818
rect -12136 13584 -12105 13818
rect -12213 13531 -12105 13584
rect -12045 13818 -11937 13871
rect -12045 13584 -12014 13818
rect -11968 13584 -11937 13818
rect -12045 13531 -11937 13584
rect -11877 13818 -11769 13871
rect -11877 13584 -11846 13818
rect -11800 13584 -11769 13818
rect -11877 13531 -11769 13584
rect -11709 13818 -11601 13871
rect -11709 13584 -11678 13818
rect -11632 13584 -11601 13818
rect -11709 13531 -11601 13584
rect -11541 13818 -11433 13871
rect -11541 13584 -11510 13818
rect -11464 13584 -11433 13818
rect -11541 13531 -11433 13584
rect -11373 13818 -11265 13871
rect -11373 13584 -11342 13818
rect -11296 13584 -11265 13818
rect -11373 13531 -11265 13584
rect -11205 13818 -11097 13871
rect -11205 13584 -11174 13818
rect -11128 13584 -11097 13818
rect -11205 13531 -11097 13584
rect -11037 13818 -10929 13871
rect -11037 13584 -11006 13818
rect -10960 13584 -10929 13818
rect -11037 13531 -10929 13584
rect -10869 13818 -10761 13871
rect -10869 13584 -10838 13818
rect -10792 13584 -10761 13818
rect -10869 13531 -10761 13584
rect -10701 13818 -10593 13871
rect -10701 13584 -10670 13818
rect -10624 13584 -10593 13818
rect -10701 13531 -10593 13584
rect -10533 13818 -10425 13871
rect -10533 13584 -10502 13818
rect -10456 13584 -10425 13818
rect -10533 13531 -10425 13584
rect -10365 13818 -10257 13871
rect -10365 13584 -10334 13818
rect -10288 13584 -10257 13818
rect -10365 13531 -10257 13584
rect -10197 13818 -10089 13871
rect -10197 13584 -10166 13818
rect -10120 13584 -10089 13818
rect -10197 13531 -10089 13584
rect -10029 13818 -9921 13871
rect -10029 13584 -9998 13818
rect -9952 13584 -9921 13818
rect -10029 13531 -9921 13584
<< ndiffc >>
rect -12710 13201 -12664 13247
rect -12542 13201 -12496 13247
rect -12374 13201 -12328 13247
rect -12206 13201 -12160 13247
rect -11930 13201 -11884 13247
rect -11762 13201 -11716 13247
rect -11594 13201 -11548 13247
rect -11426 13201 -11380 13247
rect -11258 13201 -11212 13247
rect -11090 13201 -11044 13247
rect -10922 13201 -10876 13247
rect -10754 13201 -10708 13247
rect -10478 13201 -10432 13247
rect -10310 13201 -10264 13247
rect -10142 13201 -10096 13247
rect -9974 13201 -9928 13247
<< pdiffc >>
rect -12686 13584 -12640 13818
rect -12518 13584 -12472 13818
rect -12350 13584 -12304 13818
rect -12182 13584 -12136 13818
rect -12014 13584 -11968 13818
rect -11846 13584 -11800 13818
rect -11678 13584 -11632 13818
rect -11510 13584 -11464 13818
rect -11342 13584 -11296 13818
rect -11174 13584 -11128 13818
rect -11006 13584 -10960 13818
rect -10838 13584 -10792 13818
rect -10670 13584 -10624 13818
rect -10502 13584 -10456 13818
rect -10334 13584 -10288 13818
rect -10166 13584 -10120 13818
rect -9998 13584 -9952 13818
<< psubdiff >>
rect -12594 12951 -12444 12973
rect -12594 12905 -12542 12951
rect -12496 12905 -12444 12951
rect -12594 12883 -12444 12905
rect -12354 12951 -12204 12973
rect -12354 12905 -12302 12951
rect -12256 12905 -12204 12951
rect -12354 12883 -12204 12905
rect -12114 12951 -11964 12973
rect -12114 12905 -12062 12951
rect -12016 12905 -11964 12951
rect -12114 12883 -11964 12905
rect -11874 12951 -11724 12973
rect -11874 12905 -11822 12951
rect -11776 12905 -11724 12951
rect -11874 12883 -11724 12905
rect -11634 12951 -11484 12973
rect -11634 12905 -11582 12951
rect -11536 12905 -11484 12951
rect -11634 12883 -11484 12905
rect -11394 12951 -11244 12973
rect -11394 12905 -11342 12951
rect -11296 12905 -11244 12951
rect -11394 12883 -11244 12905
rect -11154 12951 -11004 12973
rect -11154 12905 -11102 12951
rect -11056 12905 -11004 12951
rect -11154 12883 -11004 12905
rect -10914 12951 -10764 12973
rect -10914 12905 -10862 12951
rect -10816 12905 -10764 12951
rect -10914 12883 -10764 12905
rect -10674 12951 -10524 12973
rect -10674 12905 -10622 12951
rect -10576 12905 -10524 12951
rect -10674 12883 -10524 12905
rect -10434 12951 -10284 12973
rect -10434 12905 -10382 12951
rect -10336 12905 -10284 12951
rect -10434 12883 -10284 12905
rect -10194 12951 -10044 12973
rect -10194 12905 -10142 12951
rect -10096 12905 -10044 12951
rect -10194 12883 -10044 12905
<< nsubdiff >>
rect -12594 14105 -12444 14127
rect -12594 14059 -12542 14105
rect -12496 14059 -12444 14105
rect -12594 14037 -12444 14059
rect -12354 14105 -12204 14127
rect -12354 14059 -12302 14105
rect -12256 14059 -12204 14105
rect -12354 14037 -12204 14059
rect -12114 14105 -11964 14127
rect -12114 14059 -12062 14105
rect -12016 14059 -11964 14105
rect -12114 14037 -11964 14059
rect -11874 14105 -11724 14127
rect -11874 14059 -11822 14105
rect -11776 14059 -11724 14105
rect -11874 14037 -11724 14059
rect -11634 14105 -11484 14127
rect -11634 14059 -11582 14105
rect -11536 14059 -11484 14105
rect -11634 14037 -11484 14059
rect -11394 14105 -11244 14127
rect -11394 14059 -11342 14105
rect -11296 14059 -11244 14105
rect -11394 14037 -11244 14059
rect -11154 14105 -11004 14127
rect -11154 14059 -11102 14105
rect -11056 14059 -11004 14105
rect -11154 14037 -11004 14059
rect -10914 14105 -10764 14127
rect -10914 14059 -10862 14105
rect -10816 14059 -10764 14105
rect -10914 14037 -10764 14059
rect -10674 14105 -10524 14127
rect -10674 14059 -10622 14105
rect -10576 14059 -10524 14105
rect -10674 14037 -10524 14059
rect -10434 14105 -10284 14127
rect -10434 14059 -10382 14105
rect -10336 14059 -10284 14105
rect -10434 14037 -10284 14059
rect -10194 14105 -10044 14127
rect -10194 14059 -10142 14105
rect -10096 14059 -10044 14105
rect -10194 14037 -10044 14059
<< psubdiffcont >>
rect -12542 12905 -12496 12951
rect -12302 12905 -12256 12951
rect -12062 12905 -12016 12951
rect -11822 12905 -11776 12951
rect -11582 12905 -11536 12951
rect -11342 12905 -11296 12951
rect -11102 12905 -11056 12951
rect -10862 12905 -10816 12951
rect -10622 12905 -10576 12951
rect -10382 12905 -10336 12951
rect -10142 12905 -10096 12951
<< nsubdiffcont >>
rect -12542 14059 -12496 14105
rect -12302 14059 -12256 14105
rect -12062 14059 -12016 14105
rect -11822 14059 -11776 14105
rect -11582 14059 -11536 14105
rect -11342 14059 -11296 14105
rect -11102 14059 -11056 14105
rect -10862 14059 -10816 14105
rect -10622 14059 -10576 14105
rect -10382 14059 -10336 14105
rect -10142 14059 -10096 14105
<< polysilicon >>
rect -12105 13969 -10197 14009
rect -12609 13871 -12549 13921
rect -12441 13871 -12381 13921
rect -12105 13871 -12045 13969
rect -11937 13871 -11877 13921
rect -11769 13871 -11709 13921
rect -11601 13871 -11541 13921
rect -11265 13871 -11205 13969
rect -11097 13871 -11037 13921
rect -10761 13871 -10701 13921
rect -10593 13871 -10533 13921
rect -10257 13871 -10197 13969
rect -10089 13871 -10029 13921
rect -12609 13503 -12549 13531
rect -12633 13455 -12549 13503
rect -12633 13409 -12614 13455
rect -12568 13409 -12549 13455
rect -12633 13379 -12549 13409
rect -12633 13309 -12573 13379
rect -12441 13377 -12381 13531
rect -12105 13503 -12045 13531
rect -12465 13337 -12381 13377
rect -12129 13463 -12045 13503
rect -12465 13309 -12405 13337
rect -12129 13309 -12069 13463
rect -11937 13462 -11877 13531
rect -11769 13462 -11709 13531
rect -11601 13503 -11541 13531
rect -11601 13463 -11457 13503
rect -11937 13441 -11709 13462
rect -11937 13395 -11843 13441
rect -11797 13395 -11709 13441
rect -11937 13377 -11709 13395
rect -12021 13337 -11625 13377
rect -12021 13309 -11961 13337
rect -11685 13309 -11625 13337
rect -11517 13309 -11457 13463
rect -11265 13377 -11205 13531
rect -11097 13503 -11037 13531
rect -10761 13503 -10701 13531
rect -11097 13463 -10701 13503
rect -10593 13503 -10533 13531
rect -10593 13463 -10509 13503
rect -10822 13441 -10723 13463
rect -10822 13395 -10795 13441
rect -10749 13395 -10723 13441
rect -10822 13377 -10723 13395
rect -11265 13337 -11121 13377
rect -11181 13309 -11121 13337
rect -11013 13337 -10617 13377
rect -11013 13309 -10953 13337
rect -10677 13309 -10617 13337
rect -10569 13309 -10509 13463
rect -10257 13377 -10197 13531
rect -10089 13503 -10029 13531
rect -10089 13455 -10005 13503
rect -10089 13409 -10070 13455
rect -10024 13409 -10005 13455
rect -10089 13379 -10005 13409
rect -10257 13337 -10173 13377
rect -10233 13309 -10173 13337
rect -10065 13309 -10005 13379
rect -12633 13089 -12573 13139
rect -12465 13041 -12405 13139
rect -12129 13089 -12069 13139
rect -12021 13089 -11961 13139
rect -11685 13089 -11625 13139
rect -11517 13041 -11457 13139
rect -11181 13089 -11121 13139
rect -11013 13089 -10953 13139
rect -10677 13089 -10617 13139
rect -10569 13041 -10509 13139
rect -10233 13089 -10173 13139
rect -10065 13089 -10005 13139
rect -12465 13001 -10509 13041
<< polycontact >>
rect -12614 13409 -12568 13455
rect -11843 13395 -11797 13441
rect -10795 13395 -10749 13441
rect -10070 13409 -10024 13455
<< metal1 >>
rect -12624 14105 -10014 14127
rect -12624 14059 -12542 14105
rect -12496 14059 -12302 14105
rect -12256 14059 -12062 14105
rect -12016 14059 -11822 14105
rect -11776 14059 -11582 14105
rect -11536 14059 -11342 14105
rect -11296 14059 -11102 14105
rect -11056 14059 -10862 14105
rect -10816 14059 -10622 14105
rect -10576 14059 -10382 14105
rect -10336 14059 -10142 14105
rect -10096 14059 -10014 14105
rect -12624 13987 -10014 14059
rect -12690 13818 -12638 13871
rect -12690 13584 -12686 13818
rect -12640 13584 -12638 13818
rect -12690 13583 -12638 13584
rect -12743 13531 -12638 13583
rect -12521 13818 -12469 13987
rect -12521 13584 -12518 13818
rect -12472 13584 -12469 13818
rect -12521 13531 -12469 13584
rect -12354 13818 -12302 13874
rect -12354 13584 -12350 13818
rect -12304 13584 -12302 13818
rect -12743 13462 -12691 13531
rect -12354 13513 -12302 13584
rect -12185 13818 -12133 13987
rect -12185 13584 -12182 13818
rect -12136 13584 -12133 13818
rect -12185 13531 -12133 13584
rect -12017 13818 -11965 13871
rect -12017 13584 -12014 13818
rect -11968 13584 -11965 13818
rect -12792 13412 -12691 13462
rect -12792 13360 -12768 13412
rect -12716 13360 -12691 13412
rect -12633 13458 -12549 13475
rect -12633 13406 -12617 13458
rect -12565 13406 -12549 13458
rect -12633 13379 -12549 13406
rect -12378 13471 -12302 13513
rect -12378 13419 -12367 13471
rect -12315 13419 -12302 13471
rect -12792 13309 -12691 13360
rect -12378 13337 -12302 13419
rect -12743 13257 -12661 13309
rect -12713 13247 -12661 13257
rect -12713 13201 -12710 13247
rect -12664 13201 -12661 13247
rect -12713 13134 -12661 13201
rect -12545 13247 -12493 13309
rect -12545 13201 -12542 13247
rect -12496 13201 -12493 13247
rect -12545 13023 -12493 13201
rect -12378 13247 -12326 13337
rect -12017 13309 -11965 13584
rect -11849 13818 -11797 13987
rect -11849 13584 -11846 13818
rect -11800 13584 -11797 13818
rect -11849 13531 -11797 13584
rect -11681 13818 -11629 13878
rect -11681 13584 -11678 13818
rect -11632 13584 -11629 13818
rect -11681 13512 -11629 13584
rect -11541 13818 -11433 13871
rect -11541 13779 -11510 13818
rect -11464 13779 -11433 13818
rect -11541 13623 -11513 13779
rect -11461 13623 -11433 13779
rect -11541 13584 -11510 13623
rect -11464 13584 -11433 13623
rect -11541 13560 -11433 13584
rect -11345 13818 -11293 13987
rect -11345 13584 -11342 13818
rect -11296 13584 -11293 13818
rect -11345 13560 -11293 13584
rect -11177 13818 -11125 13871
rect -11177 13584 -11174 13818
rect -11128 13584 -11125 13818
rect -11177 13512 -11125 13584
rect -11037 13818 -10929 13871
rect -11037 13779 -11006 13818
rect -10960 13779 -10929 13818
rect -11037 13623 -11009 13779
rect -10957 13623 -10929 13779
rect -11037 13584 -11006 13623
rect -10960 13584 -10929 13623
rect -11037 13560 -10929 13584
rect -10841 13818 -10789 13987
rect -10841 13584 -10838 13818
rect -10792 13584 -10789 13818
rect -10841 13531 -10789 13584
rect -10673 13818 -10621 13871
rect -10673 13584 -10670 13818
rect -10624 13584 -10621 13818
rect -11902 13444 -11745 13462
rect -11681 13460 -11125 13512
rect -11902 13392 -11846 13444
rect -11794 13392 -11745 13444
rect -10822 13444 -10723 13463
rect -11902 13377 -11745 13392
rect -11429 13357 -10873 13409
rect -10822 13392 -10798 13444
rect -10746 13392 -10723 13444
rect -10822 13377 -10723 13392
rect -12378 13201 -12374 13247
rect -12328 13201 -12326 13247
rect -12378 13139 -12326 13201
rect -12209 13247 -12157 13309
rect -12209 13201 -12206 13247
rect -12160 13201 -12157 13247
rect -12209 13023 -12157 13201
rect -12021 13249 -11853 13309
rect -12021 13197 -12006 13249
rect -11954 13247 -11853 13249
rect -11954 13201 -11930 13247
rect -11884 13201 -11853 13247
rect -11954 13197 -11853 13201
rect -12021 13139 -11853 13197
rect -11766 13247 -11714 13309
rect -11766 13201 -11762 13247
rect -11716 13201 -11714 13247
rect -11766 13123 -11714 13201
rect -11625 13251 -11517 13285
rect -11625 13199 -11597 13251
rect -11545 13199 -11517 13251
rect -11625 13171 -11517 13199
rect -11429 13247 -11377 13357
rect -11429 13201 -11426 13247
rect -11380 13201 -11377 13247
rect -11429 13171 -11377 13201
rect -11261 13247 -11209 13309
rect -11261 13201 -11258 13247
rect -11212 13201 -11209 13247
rect -11261 13123 -11209 13201
rect -11766 13071 -11209 13123
rect -11094 13247 -11042 13309
rect -11094 13201 -11090 13247
rect -11044 13201 -11042 13247
rect -11094 13023 -11042 13201
rect -10925 13247 -10873 13357
rect -10673 13309 -10621 13584
rect -10505 13818 -10453 13987
rect -10505 13584 -10502 13818
rect -10456 13584 -10453 13818
rect -10505 13531 -10453 13584
rect -10337 13818 -10285 13874
rect -10337 13584 -10334 13818
rect -10288 13584 -10285 13818
rect -10337 13513 -10285 13584
rect -10169 13818 -10117 13987
rect -10169 13584 -10166 13818
rect -10120 13584 -10117 13818
rect -10169 13531 -10117 13584
rect -10001 13818 -9949 13871
rect -10001 13584 -9998 13818
rect -9952 13584 -9949 13818
rect -10001 13583 -9949 13584
rect -10001 13531 -9897 13583
rect -10337 13471 -10261 13513
rect -10337 13419 -10324 13471
rect -10272 13419 -10261 13471
rect -10337 13377 -10261 13419
rect -10089 13458 -10005 13480
rect -10089 13406 -10073 13458
rect -10021 13406 -10005 13458
rect -10089 13379 -10005 13406
rect -9949 13462 -9897 13531
rect -9949 13412 -9846 13462
rect -10925 13201 -10922 13247
rect -10876 13201 -10873 13247
rect -10925 13139 -10873 13201
rect -10785 13249 -10617 13309
rect -10785 13247 -10691 13249
rect -10785 13201 -10754 13247
rect -10708 13201 -10691 13247
rect -10785 13197 -10691 13201
rect -10639 13197 -10617 13249
rect -10785 13139 -10617 13197
rect -10481 13247 -10429 13309
rect -10481 13201 -10478 13247
rect -10432 13201 -10429 13247
rect -10481 13023 -10429 13201
rect -10313 13247 -10261 13377
rect -9949 13360 -9921 13412
rect -9869 13360 -9846 13412
rect -9949 13309 -9846 13360
rect -10313 13201 -10310 13247
rect -10264 13201 -10261 13247
rect -10313 13139 -10261 13201
rect -10145 13247 -10093 13309
rect -10145 13201 -10142 13247
rect -10096 13201 -10093 13247
rect -10145 13023 -10093 13201
rect -9977 13257 -9897 13309
rect -9977 13247 -9925 13257
rect -9977 13201 -9974 13247
rect -9928 13201 -9925 13247
rect -9977 13140 -9925 13201
rect -12624 12951 -10014 13023
rect -12624 12905 -12542 12951
rect -12496 12905 -12302 12951
rect -12256 12905 -12062 12951
rect -12016 12905 -11822 12951
rect -11776 12905 -11582 12951
rect -11536 12905 -11342 12951
rect -11296 12905 -11102 12951
rect -11056 12905 -10862 12951
rect -10816 12905 -10622 12951
rect -10576 12905 -10382 12951
rect -10336 12905 -10142 12951
rect -10096 12905 -10014 12951
rect -12624 12883 -10014 12905
<< via1 >>
rect -12768 13360 -12716 13412
rect -12617 13455 -12565 13458
rect -12617 13409 -12614 13455
rect -12614 13409 -12568 13455
rect -12568 13409 -12565 13455
rect -12617 13406 -12565 13409
rect -12367 13419 -12315 13471
rect -11513 13623 -11510 13779
rect -11510 13623 -11464 13779
rect -11464 13623 -11461 13779
rect -11009 13623 -11006 13779
rect -11006 13623 -10960 13779
rect -10960 13623 -10957 13779
rect -11846 13441 -11794 13444
rect -11846 13395 -11843 13441
rect -11843 13395 -11797 13441
rect -11797 13395 -11794 13441
rect -11846 13392 -11794 13395
rect -10798 13441 -10746 13444
rect -10798 13395 -10795 13441
rect -10795 13395 -10749 13441
rect -10749 13395 -10746 13441
rect -10798 13392 -10746 13395
rect -12006 13197 -11954 13249
rect -11597 13247 -11545 13251
rect -11597 13201 -11594 13247
rect -11594 13201 -11548 13247
rect -11548 13201 -11545 13247
rect -11597 13199 -11545 13201
rect -10324 13419 -10272 13471
rect -10073 13455 -10021 13458
rect -10073 13409 -10070 13455
rect -10070 13409 -10024 13455
rect -10024 13409 -10021 13455
rect -10073 13406 -10021 13409
rect -10691 13197 -10639 13249
rect -9921 13360 -9869 13412
<< metal2 >>
rect -11601 13779 -11433 13871
rect -11601 13623 -11513 13779
rect -11461 13730 -11433 13779
rect -11037 13779 -10929 13871
rect -11037 13730 -11009 13779
rect -11461 13670 -11009 13730
rect -11461 13623 -11433 13670
rect -11601 13560 -11433 13623
rect -11037 13623 -11009 13670
rect -10957 13623 -10929 13779
rect -11037 13560 -10929 13623
rect -12633 13475 -12573 13503
rect -12792 13412 -12693 13462
rect -12792 13360 -12768 13412
rect -12716 13360 -12693 13412
rect -12792 13309 -12693 13360
rect -12633 13458 -12549 13475
rect -12633 13406 -12617 13458
rect -12565 13406 -12549 13458
rect -12633 13379 -12549 13406
rect -12378 13471 -12302 13513
rect -12378 13419 -12367 13471
rect -12315 13450 -12302 13471
rect -11937 13450 -11709 13462
rect -12315 13444 -11709 13450
rect -12315 13419 -11846 13444
rect -12378 13392 -11846 13419
rect -11794 13392 -11709 13444
rect -12378 13390 -11709 13392
rect -12633 13199 -12573 13379
rect -12378 13337 -12302 13390
rect -11937 13377 -11709 13390
rect -12021 13249 -11853 13309
rect -11601 13285 -11541 13560
rect -10337 13471 -10261 13513
rect -10065 13480 -10005 13503
rect -10822 13444 -10723 13463
rect -10822 13392 -10798 13444
rect -10746 13437 -10723 13444
rect -10337 13437 -10324 13471
rect -10746 13419 -10324 13437
rect -10272 13419 -10261 13471
rect -10746 13392 -10261 13419
rect -10822 13377 -10261 13392
rect -10089 13458 -10005 13480
rect -10089 13406 -10073 13458
rect -10021 13406 -10005 13458
rect -10089 13379 -10005 13406
rect -12021 13199 -12006 13249
rect -12633 13197 -12006 13199
rect -11954 13197 -11853 13249
rect -12633 13139 -11853 13197
rect -11625 13251 -11517 13285
rect -11625 13199 -11597 13251
rect -11545 13199 -11517 13251
rect -11625 13171 -11517 13199
rect -10785 13249 -10617 13309
rect -10785 13197 -10691 13249
rect -10639 13199 -10617 13249
rect -10065 13199 -10005 13379
rect -9945 13412 -9846 13462
rect -9945 13360 -9921 13412
rect -9869 13360 -9846 13412
rect -9945 13309 -9846 13360
rect -10639 13197 -10005 13199
rect -11601 13152 -11541 13171
rect -10785 13139 -10005 13197
<< labels >>
flabel metal2 s -12768 13343 -12768 13343 2 FreeSans 560 0 0 0 L
port 1 nsew
flabel metal2 s -11586 13378 -11586 13378 2 FreeSans 560 0 0 0 E
port 2 nsew
flabel metal2 s -9881 13336 -9881 13336 2 FreeSans 560 0 0 0 G
port 3 nsew
flabel metal1 s -10244 14085 -10244 14085 2 FreeSans 460 0 0 0 VDD
port 4 nsew
flabel metal1 s -10244 12936 -10244 12936 2 FreeSans 460 0 0 0 VSS
port 5 nsew
rlabel polysilicon s -12410 13400 -12410 13400 4 A
port 7 se
rlabel polysilicon s -12070 13910 -12070 13910 4 B
port 6 se
<< end >>
