* NGSPICE file created from 2bit_comp_1x.ext - technology: gf180mcuD

.subckt x2bit_comp_1x VDD VSS B0 A0 B1 A1 L G E
X0 my_xor_0.Y a_700_n970# a_600_n920# VDD pfet_03v3 ad=0.7225p pd=2.55u as=0.425p ps=2.2u w=1.7u l=0.3u
X1 a_2910_n920# E G VDD pfet_03v3 ad=0.935p pd=4.5u as=0.4675p ps=2.25u w=1.7u l=0.3u
X2 VDD my_nxor_0.Y a_1240_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.935p ps=4.5u w=1.7u l=0.3u
X3 my_nand_0.Y my_nxor_0.Y a_1880_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
X4 VSS a_3100_610# a_3390_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2125p ps=1.35u w=0.85u l=0.3u
X5 VDD my_nand_0.B my_nand_0.Y VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X6 a_3390_720# a_2670_210# L VDD pfet_03v3 ad=0.425p pd=2.2u as=0.7225p ps=2.55u w=1.7u l=0.3u
X7 a_3000_210# my_nor_0.Y VSS VSS nfet_03v3 ad=0.2125p pd=1.35u as=0.23375p ps=1.4u w=0.85u l=0.3u
X8 VDD my_xor_0.Y my_nand_0.B VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X9 VDD my_nor_0.Y a_2670_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X10 VSS a_700_n970# a_990_n240# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2125p ps=1.35u w=0.85u l=0.3u
X11 a_3250_n920# L VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.4675p ps=2.25u w=1.7u l=0.3u
X12 a_990_n240# a_270_n920# my_xor_0.Y VSS nfet_03v3 ad=0.2125p pd=1.35u as=0.36125p ps=1.7u w=0.85u l=0.3u
X13 a_1580_720# my_nxor_0.Y VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.4675p ps=2.25u w=1.7u l=0.3u
X14 a_2460_n920# my_nand_0.Y VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.4675p ps=2.25u w=1.7u l=0.3u
X15 VDD my_nand_0.Y a_3390_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.425p ps=2.2u w=1.7u l=0.3u
X16 a_3100_610# my_nand_0.Y VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X17 a_3000_720# my_nor_0.Y VDD VDD pfet_03v3 ad=0.425p pd=2.2u as=0.4675p ps=2.25u w=1.7u l=0.3u
X18 L my_nand_0.Y a_3000_210# VSS nfet_03v3 ad=0.36125p pd=1.7u as=0.2125p ps=1.35u w=0.85u l=0.3u
X19 VSS A1 a_780_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.14875p ps=1.2u w=0.85u l=0.3u
X20 a_1820_n240# B0 my_nand_0.B VSS nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
X21 VSS my_xor_0.Y E VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X22 a_600_n920# B0 VDD VDD pfet_03v3 ad=0.425p pd=2.2u as=0.4675p ps=2.25u w=1.7u l=0.3u
X23 a_2120_n920# my_xor_0.Y E VDD pfet_03v3 ad=0.935p pd=4.5u as=0.4675p ps=2.25u w=1.7u l=0.3u
X24 VSS B1 a_90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X25 a_780_210# a_90_210# my_nxor_0.Y VSS nfet_03v3 ad=0.14875p pd=1.2u as=0.37375p ps=1.75u w=0.85u l=0.3u
X26 G E a_3250_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X27 a_3100_610# my_nand_0.Y VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X28 VSS my_nand_0.B a_2220_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.10625p ps=1.1u w=0.85u l=0.3u
X29 VSS B0 a_270_n920# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X30 VDD A1 a_780_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.2975p ps=2.05u w=1.7u l=0.3u
X31 L a_3100_610# a_3000_720# VDD pfet_03v3 ad=0.7225p pd=2.55u as=0.425p ps=2.2u w=1.7u l=0.3u
X32 my_nxor_0.Y a_490_160# a_420_210# VSS nfet_03v3 ad=0.37375p pd=1.75u as=0.14875p ps=1.2u w=0.85u l=0.3u
X33 VDD L a_2910_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.935p ps=4.5u w=1.7u l=0.3u
X34 VDD B1 a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X35 a_780_720# B1 my_nxor_0.Y VDD pfet_03v3 ad=0.2975p pd=2.05u as=0.7225p ps=2.55u w=1.7u l=0.3u
X36 a_420_210# B1 VSS VSS nfet_03v3 ad=0.14875p pd=1.2u as=0.23375p ps=1.4u w=0.85u l=0.3u
X37 a_700_n970# A0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X38 a_1480_n240# my_xor_0.Y VSS VSS nfet_03v3 ad=0.4675p pd=2.8u as=0.23375p ps=1.4u w=0.85u l=0.3u
X39 a_490_160# A1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X40 my_nor_0.Y my_nxor_0.Y VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X41 my_xor_0.Y A0 a_600_n240# VSS nfet_03v3 ad=0.36125p pd=1.7u as=0.2125p ps=1.35u w=0.85u l=0.3u
X42 a_1880_210# my_nand_0.B VSS VSS nfet_03v3 ad=0.4675p pd=2.8u as=0.23375p ps=1.4u w=0.85u l=0.3u
X43 G L VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X44 VDD A0 a_990_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.425p ps=2.2u w=1.7u l=0.3u
X45 my_nxor_0.Y a_490_160# a_420_720# VDD pfet_03v3 ad=0.7225p pd=2.55u as=0.2975p ps=2.05u w=1.7u l=0.3u
X46 a_990_n920# a_270_n920# my_xor_0.Y VDD pfet_03v3 ad=0.425p pd=2.2u as=0.7225p ps=2.55u w=1.7u l=0.3u
X47 my_nor_0.Y B1 a_1580_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X48 my_nand_0.B B0 VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X49 E my_xor_0.Y a_2460_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X50 a_420_720# a_90_210# VDD VDD pfet_03v3 ad=0.2975p pd=2.05u as=0.4675p ps=2.25u w=1.7u l=0.3u
X51 a_490_160# A1 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X52 VSS B1 my_nor_0.Y VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X53 VSS my_xor_0.Y a_1820_n240# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.10625p ps=1.1u w=0.85u l=0.3u
X54 VDD my_nand_0.Y a_2120_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.935p ps=4.5u w=1.7u l=0.3u
X55 a_1240_720# B1 my_nor_0.Y VDD pfet_03v3 ad=0.935p pd=4.5u as=0.4675p ps=2.25u w=1.7u l=0.3u
X56 a_600_n240# B0 VSS VSS nfet_03v3 ad=0.2125p pd=1.35u as=0.23375p ps=1.4u w=0.85u l=0.3u
X57 a_3390_210# a_2670_210# L VSS nfet_03v3 ad=0.2125p pd=1.35u as=0.36125p ps=1.7u w=0.85u l=0.3u
X58 my_nand_0.B B0 a_1480_n240# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
X59 E my_nand_0.Y VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X60 VDD B0 a_270_n920# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X61 my_nand_0.Y my_nxor_0.Y VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X62 VSS my_nor_0.Y a_2670_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X63 a_2220_210# my_nxor_0.Y my_nand_0.Y VSS nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
X64 VSS E G VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X65 a_700_n970# A0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
.ends

