magic
tech gf180mcuD
timestamp 1755257261
<< nwell >>
rect 0 63 387 127
rect 30 -113 347 -49
<< nmos >>
rect 19 21 25 38
rect 36 21 42 38
rect 49 21 55 38
rect 72 21 78 38
rect 85 21 91 38
rect 102 21 108 38
rect 147 21 153 38
rect 164 21 170 38
rect 213 21 219 38
rect 224 21 230 38
rect 272 21 278 38
rect 289 21 295 38
rect 305 21 311 38
rect 328 21 334 38
rect 344 21 350 38
rect 361 21 367 38
rect 49 -24 55 -7
rect 66 -24 72 -7
rect 82 -24 88 -7
rect 105 -24 111 -7
rect 121 -24 127 -7
rect 138 -24 144 -7
rect 180 -24 186 -7
rect 191 -24 197 -7
rect 240 -24 246 -7
rect 257 -24 263 -7
rect 302 -24 308 -7
rect 319 -24 325 -7
<< pmos >>
rect 19 72 25 106
rect 36 72 42 106
rect 49 72 55 106
rect 72 72 78 106
rect 85 72 91 106
rect 102 72 108 106
rect 150 72 156 106
rect 161 72 167 106
rect 210 72 216 106
rect 227 72 233 106
rect 272 72 278 106
rect 289 72 295 106
rect 305 72 311 106
rect 328 72 334 106
rect 344 72 350 106
rect 361 72 367 106
rect 49 -92 55 -58
rect 66 -92 72 -58
rect 82 -92 88 -58
rect 105 -92 111 -58
rect 121 -92 127 -58
rect 138 -92 144 -58
rect 177 -92 183 -58
rect 194 -92 200 -58
rect 243 -92 249 -58
rect 254 -92 260 -58
rect 305 -92 311 -58
rect 316 -92 322 -58
<< ndiff >>
rect 58 38 68 39
rect 9 36 19 38
rect 9 23 11 36
rect 16 23 19 36
rect 9 21 19 23
rect 25 36 36 38
rect 25 23 28 36
rect 33 23 36 36
rect 25 21 36 23
rect 42 21 49 38
rect 55 37 72 38
rect 55 23 61 37
rect 66 23 72 37
rect 55 21 72 23
rect 78 21 85 38
rect 91 36 102 38
rect 91 23 94 36
rect 99 23 102 36
rect 91 21 102 23
rect 108 36 118 38
rect 108 23 111 36
rect 116 23 118 36
rect 108 21 118 23
rect 137 36 147 38
rect 137 23 139 36
rect 144 23 147 36
rect 137 21 147 23
rect 153 36 164 38
rect 153 23 156 36
rect 161 23 164 36
rect 153 21 164 23
rect 170 36 180 38
rect 170 23 173 36
rect 178 23 180 36
rect 170 21 180 23
rect 203 29 213 38
rect 203 23 205 29
rect 210 23 213 29
rect 203 21 213 23
rect 219 21 224 38
rect 230 36 240 38
rect 230 23 233 36
rect 238 23 240 36
rect 230 21 240 23
rect 262 36 272 38
rect 262 23 264 36
rect 269 23 272 36
rect 262 21 272 23
rect 278 36 289 38
rect 278 23 281 36
rect 286 23 289 36
rect 278 21 289 23
rect 295 21 305 38
rect 311 28 328 38
rect 311 23 317 28
rect 322 23 328 28
rect 311 21 328 23
rect 334 21 344 38
rect 350 35 361 38
rect 350 23 353 35
rect 358 23 361 35
rect 350 21 361 23
rect 367 36 377 38
rect 367 23 370 36
rect 375 23 377 36
rect 367 21 377 23
rect 39 -9 49 -7
rect 39 -22 41 -9
rect 46 -22 49 -9
rect 39 -24 49 -22
rect 55 -9 66 -7
rect 55 -22 58 -9
rect 63 -22 66 -9
rect 55 -24 66 -22
rect 72 -24 82 -7
rect 88 -9 105 -7
rect 88 -14 94 -9
rect 99 -14 105 -9
rect 88 -24 105 -14
rect 111 -24 121 -7
rect 127 -9 138 -7
rect 127 -21 130 -9
rect 135 -21 138 -9
rect 127 -24 138 -21
rect 144 -9 154 -7
rect 144 -22 147 -9
rect 152 -22 154 -9
rect 144 -24 154 -22
rect 170 -9 180 -7
rect 170 -15 172 -9
rect 177 -15 180 -9
rect 170 -24 180 -15
rect 186 -24 191 -7
rect 197 -9 207 -7
rect 197 -22 200 -9
rect 205 -22 207 -9
rect 197 -24 207 -22
rect 230 -9 240 -7
rect 230 -22 232 -9
rect 237 -22 240 -9
rect 230 -24 240 -22
rect 246 -9 257 -7
rect 246 -22 249 -9
rect 254 -22 257 -9
rect 246 -24 257 -22
rect 263 -9 273 -7
rect 263 -22 266 -9
rect 271 -22 273 -9
rect 263 -24 273 -22
rect 292 -9 302 -7
rect 292 -22 294 -9
rect 299 -22 302 -9
rect 292 -24 302 -22
rect 308 -9 319 -7
rect 308 -22 311 -9
rect 316 -22 319 -9
rect 308 -24 319 -22
rect 325 -9 335 -7
rect 325 -22 328 -9
rect 333 -22 335 -9
rect 325 -24 335 -22
<< pdiff >>
rect 9 104 19 106
rect 9 96 11 104
rect 16 96 19 104
rect 9 72 19 96
rect 25 104 36 106
rect 25 96 28 104
rect 33 96 36 104
rect 25 72 36 96
rect 42 72 49 106
rect 55 104 72 106
rect 55 96 61 104
rect 66 96 72 104
rect 55 72 72 96
rect 78 72 85 106
rect 91 104 102 106
rect 91 96 94 104
rect 99 96 102 104
rect 91 72 102 96
rect 108 104 118 106
rect 108 96 111 104
rect 116 96 118 104
rect 108 72 118 96
rect 140 104 150 106
rect 140 74 142 104
rect 147 74 150 104
rect 140 72 150 74
rect 156 72 161 106
rect 167 104 177 106
rect 167 81 170 104
rect 175 81 177 104
rect 167 72 177 81
rect 200 104 210 106
rect 200 74 202 104
rect 207 74 210 104
rect 200 72 210 74
rect 216 104 227 106
rect 216 79 219 104
rect 224 79 227 104
rect 216 72 227 79
rect 233 104 243 106
rect 233 74 236 104
rect 241 74 243 104
rect 233 72 243 74
rect 262 104 272 106
rect 262 74 264 104
rect 269 74 272 104
rect 262 72 272 74
rect 278 104 289 106
rect 278 80 281 104
rect 286 80 289 104
rect 278 72 289 80
rect 295 72 305 106
rect 311 104 328 106
rect 311 99 317 104
rect 322 99 328 104
rect 311 72 328 99
rect 334 72 344 106
rect 350 104 361 106
rect 350 80 353 104
rect 358 80 361 104
rect 350 72 361 80
rect 367 104 377 106
rect 367 74 370 104
rect 375 74 377 104
rect 367 72 377 74
rect 39 -60 49 -58
rect 39 -90 41 -60
rect 46 -90 49 -60
rect 39 -92 49 -90
rect 55 -66 66 -58
rect 55 -90 58 -66
rect 63 -90 66 -66
rect 55 -92 66 -90
rect 72 -92 82 -58
rect 88 -85 105 -58
rect 88 -90 94 -85
rect 99 -90 105 -85
rect 88 -92 105 -90
rect 111 -92 121 -58
rect 127 -66 138 -58
rect 127 -90 130 -66
rect 135 -90 138 -66
rect 127 -92 138 -90
rect 144 -60 154 -58
rect 144 -90 147 -60
rect 152 -90 154 -60
rect 144 -92 154 -90
rect 167 -60 177 -58
rect 167 -90 169 -60
rect 174 -90 177 -60
rect 167 -92 177 -90
rect 183 -65 194 -58
rect 183 -90 186 -65
rect 191 -90 194 -65
rect 183 -92 194 -90
rect 200 -60 210 -58
rect 200 -90 203 -60
rect 208 -90 210 -60
rect 200 -92 210 -90
rect 233 -60 243 -58
rect 233 -90 235 -60
rect 240 -90 243 -60
rect 233 -92 243 -90
rect 249 -92 254 -58
rect 260 -67 270 -58
rect 260 -90 263 -67
rect 268 -90 270 -67
rect 260 -92 270 -90
rect 295 -60 305 -58
rect 295 -90 297 -60
rect 302 -90 305 -60
rect 295 -92 305 -90
rect 311 -92 316 -58
rect 322 -67 332 -58
rect 322 -90 325 -67
rect 330 -90 332 -67
rect 322 -92 332 -90
<< ndiffc >>
rect 11 23 16 36
rect 28 23 33 36
rect 61 23 66 37
rect 94 23 99 36
rect 111 23 116 36
rect 139 23 144 36
rect 156 23 161 36
rect 173 23 178 36
rect 205 23 210 29
rect 233 23 238 36
rect 264 23 269 36
rect 281 23 286 36
rect 317 23 322 28
rect 353 23 358 35
rect 370 23 375 36
rect 41 -22 46 -9
rect 58 -22 63 -9
rect 94 -14 99 -9
rect 130 -21 135 -9
rect 147 -22 152 -9
rect 172 -15 177 -9
rect 200 -22 205 -9
rect 232 -22 237 -9
rect 249 -22 254 -9
rect 266 -22 271 -9
rect 294 -22 299 -9
rect 311 -22 316 -9
rect 328 -22 333 -9
<< pdiffc >>
rect 11 96 16 104
rect 28 96 33 104
rect 61 96 66 104
rect 94 96 99 104
rect 111 96 116 104
rect 142 74 147 104
rect 170 81 175 104
rect 202 74 207 104
rect 219 79 224 104
rect 236 74 241 104
rect 264 74 269 104
rect 281 80 286 104
rect 317 99 322 104
rect 353 80 358 104
rect 370 74 375 104
rect 41 -90 46 -60
rect 58 -90 63 -66
rect 94 -90 99 -85
rect 130 -90 135 -66
rect 147 -90 152 -60
rect 169 -90 174 -60
rect 186 -90 191 -65
rect 203 -90 208 -60
rect 235 -90 240 -60
rect 263 -90 268 -67
rect 297 -90 302 -60
rect 325 -90 330 -67
<< psubdiff >>
rect 6 12 21 14
rect 6 2 11 12
rect 16 2 21 12
rect 6 0 21 2
rect 30 12 45 14
rect 30 2 35 12
rect 40 2 45 12
rect 30 0 45 2
rect 54 12 69 14
rect 54 2 59 12
rect 64 2 69 12
rect 54 0 69 2
rect 78 12 93 14
rect 78 2 83 12
rect 88 2 93 12
rect 78 0 93 2
rect 102 12 117 14
rect 102 2 107 12
rect 112 2 117 12
rect 102 0 117 2
rect 134 12 149 14
rect 134 2 139 12
rect 144 2 149 12
rect 134 0 149 2
rect 158 12 173 14
rect 158 2 163 12
rect 168 2 173 12
rect 158 0 173 2
rect 197 12 212 14
rect 197 2 202 12
rect 207 2 212 12
rect 197 0 212 2
rect 221 12 236 14
rect 221 2 226 12
rect 231 2 236 12
rect 221 0 236 2
rect 259 12 274 14
rect 259 2 264 12
rect 269 2 274 12
rect 259 0 274 2
rect 283 12 298 14
rect 283 2 288 12
rect 293 2 298 12
rect 307 12 322 14
rect 307 7 312 12
rect 317 7 322 12
rect 307 5 322 7
rect 331 12 346 14
rect 331 7 336 12
rect 341 7 346 12
rect 331 5 346 7
rect 355 12 370 14
rect 355 7 360 12
rect 365 7 370 12
rect 355 5 370 7
rect 283 0 298 2
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
rect 54 120 69 122
rect 54 115 59 120
rect 64 115 69 120
rect 54 113 69 115
rect 78 120 93 122
rect 78 115 83 120
rect 88 115 93 120
rect 78 113 93 115
rect 102 120 117 122
rect 102 115 107 120
rect 112 115 117 120
rect 102 113 117 115
rect 134 120 149 122
rect 134 115 139 120
rect 144 115 149 120
rect 134 113 149 115
rect 158 120 173 122
rect 158 115 163 120
rect 168 115 173 120
rect 158 113 173 115
rect 197 120 212 122
rect 197 115 202 120
rect 207 115 212 120
rect 197 113 212 115
rect 221 120 236 122
rect 221 115 226 120
rect 231 115 236 120
rect 221 113 236 115
rect 259 120 274 122
rect 259 115 264 120
rect 269 115 274 120
rect 259 113 274 115
rect 283 120 298 122
rect 283 115 288 120
rect 293 115 298 120
rect 283 113 298 115
rect 307 120 322 122
rect 307 115 312 120
rect 317 115 322 120
rect 307 113 322 115
rect 331 120 346 122
rect 331 115 336 120
rect 341 115 346 120
rect 331 113 346 115
rect 355 120 370 122
rect 355 115 360 120
rect 365 115 370 120
rect 355 113 370 115
rect 36 -101 51 -99
rect 36 -106 41 -101
rect 46 -106 51 -101
rect 36 -108 51 -106
rect 60 -101 75 -99
rect 60 -106 65 -101
rect 70 -106 75 -101
rect 60 -108 75 -106
rect 84 -101 99 -99
rect 84 -106 89 -101
rect 94 -106 99 -101
rect 84 -108 99 -106
rect 108 -101 123 -99
rect 108 -106 113 -101
rect 118 -106 123 -101
rect 108 -108 123 -106
rect 132 -101 147 -99
rect 132 -106 137 -101
rect 142 -106 147 -101
rect 132 -108 147 -106
rect 164 -101 179 -99
rect 164 -106 169 -101
rect 174 -106 179 -101
rect 164 -108 179 -106
rect 188 -101 203 -99
rect 188 -106 193 -101
rect 198 -106 203 -101
rect 188 -108 203 -106
rect 227 -101 242 -99
rect 227 -106 232 -101
rect 237 -106 242 -101
rect 227 -108 242 -106
rect 251 -101 266 -99
rect 251 -106 256 -101
rect 261 -106 266 -101
rect 251 -108 266 -106
rect 289 -101 304 -99
rect 289 -106 294 -101
rect 299 -106 304 -101
rect 289 -108 304 -106
rect 313 -101 328 -99
rect 313 -106 318 -101
rect 323 -106 328 -101
rect 313 -108 328 -106
<< psubdiffcont >>
rect 11 2 16 12
rect 35 2 40 12
rect 59 2 64 12
rect 83 2 88 12
rect 107 2 112 12
rect 139 2 144 12
rect 163 2 168 12
rect 202 2 207 12
rect 226 2 231 12
rect 264 2 269 12
rect 288 2 293 12
rect 312 7 317 12
rect 336 7 341 12
rect 360 7 365 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
rect 59 115 64 120
rect 83 115 88 120
rect 107 115 112 120
rect 139 115 144 120
rect 163 115 168 120
rect 202 115 207 120
rect 226 115 231 120
rect 264 115 269 120
rect 288 115 293 120
rect 312 115 317 120
rect 336 115 341 120
rect 360 115 365 120
rect 41 -106 46 -101
rect 65 -106 70 -101
rect 89 -106 94 -101
rect 113 -106 118 -101
rect 137 -106 142 -101
rect 169 -106 174 -101
rect 193 -106 198 -101
rect 232 -106 237 -101
rect 256 -106 261 -101
rect 294 -106 299 -101
rect 318 -106 323 -101
<< polysilicon >>
rect 19 106 25 111
rect 36 106 42 111
rect 49 106 55 111
rect 72 106 78 111
rect 85 106 91 111
rect 102 106 108 111
rect 150 106 156 111
rect 161 106 167 111
rect 210 106 216 111
rect 227 106 233 111
rect 272 106 278 111
rect 289 106 295 111
rect 305 106 311 111
rect 328 106 334 111
rect 344 106 350 111
rect 361 106 367 111
rect 19 54 25 72
rect 36 70 42 72
rect 31 68 42 70
rect 31 62 33 68
rect 39 62 42 68
rect 31 60 42 62
rect 49 70 55 72
rect 72 70 78 72
rect 85 70 91 72
rect 102 70 108 72
rect 49 68 63 70
rect 49 62 55 68
rect 61 62 63 68
rect 49 60 63 62
rect 70 68 80 70
rect 70 62 72 68
rect 78 62 80 68
rect 85 65 108 70
rect 150 68 156 72
rect 70 60 80 62
rect 19 52 35 54
rect 19 46 27 52
rect 33 51 35 52
rect 33 46 42 51
rect 19 44 42 46
rect 19 38 25 44
rect 36 38 42 44
rect 49 38 55 60
rect 102 54 108 65
rect 147 63 156 68
rect 161 69 167 72
rect 161 67 170 69
rect 161 65 178 67
rect 161 63 170 65
rect 147 54 153 63
rect 60 52 70 54
rect 91 52 108 54
rect 60 46 62 52
rect 68 46 78 52
rect 91 49 93 52
rect 60 44 78 46
rect 72 38 78 44
rect 85 46 93 49
rect 99 46 108 52
rect 85 44 108 46
rect 139 52 153 54
rect 139 46 142 52
rect 148 46 153 52
rect 139 44 153 46
rect 85 38 91 44
rect 102 38 108 44
rect 147 38 153 44
rect 164 59 170 63
rect 176 59 178 65
rect 164 57 178 59
rect 164 38 170 57
rect 210 54 216 72
rect 202 52 216 54
rect 202 46 205 52
rect 211 46 216 52
rect 202 44 216 46
rect 210 43 216 44
rect 227 67 233 72
rect 272 70 278 72
rect 289 70 295 72
rect 227 65 241 67
rect 227 59 233 65
rect 239 59 241 65
rect 227 57 241 59
rect 272 65 295 70
rect 305 70 311 72
rect 328 70 334 72
rect 305 68 315 70
rect 227 43 233 57
rect 210 40 219 43
rect 213 38 219 40
rect 224 40 233 43
rect 272 54 278 65
rect 305 63 307 68
rect 313 63 315 68
rect 305 61 315 63
rect 324 68 334 70
rect 324 62 326 68
rect 332 62 334 68
rect 344 70 350 72
rect 361 70 367 72
rect 344 65 367 70
rect 324 60 334 62
rect 272 52 285 54
rect 272 46 277 52
rect 283 46 285 52
rect 272 44 285 46
rect 300 48 311 50
rect 272 40 295 44
rect 300 42 302 48
rect 308 42 311 48
rect 300 40 311 42
rect 224 38 230 40
rect 272 38 278 40
rect 289 38 295 40
rect 305 38 311 40
rect 328 38 334 60
rect 340 58 350 60
rect 340 53 342 58
rect 348 53 350 58
rect 361 54 367 65
rect 340 51 350 53
rect 344 38 350 51
rect 355 52 367 54
rect 355 46 357 52
rect 363 46 367 52
rect 355 44 367 46
rect 361 38 367 44
rect 19 16 25 21
rect 36 16 42 21
rect 49 16 55 21
rect 72 16 78 21
rect 85 16 91 21
rect 102 16 108 21
rect 147 16 153 21
rect 164 16 170 21
rect 213 16 219 21
rect 224 16 230 21
rect 272 16 278 21
rect 289 16 295 21
rect 305 16 311 21
rect 328 16 334 21
rect 344 16 350 21
rect 361 16 367 21
rect 49 -7 55 -2
rect 66 -7 72 -2
rect 82 -7 88 -2
rect 105 -7 111 -2
rect 121 -7 127 -2
rect 138 -7 144 -2
rect 180 -7 186 -2
rect 191 -7 197 -2
rect 240 -7 246 -2
rect 257 -7 263 -2
rect 302 -7 308 -2
rect 319 -7 325 -2
rect 49 -26 55 -24
rect 66 -26 72 -24
rect 82 -26 88 -24
rect 49 -30 72 -26
rect 77 -28 88 -26
rect 49 -32 62 -30
rect 49 -38 54 -32
rect 60 -38 62 -32
rect 77 -34 79 -28
rect 85 -34 88 -28
rect 77 -36 88 -34
rect 49 -40 62 -38
rect 49 -51 55 -40
rect 105 -46 111 -24
rect 121 -37 127 -24
rect 138 -30 144 -24
rect 180 -26 186 -24
rect 177 -29 186 -26
rect 191 -26 197 -24
rect 191 -29 200 -26
rect 177 -30 183 -29
rect 117 -39 127 -37
rect 117 -44 119 -39
rect 125 -44 127 -39
rect 132 -32 144 -30
rect 132 -38 134 -32
rect 140 -38 144 -32
rect 132 -40 144 -38
rect 169 -32 183 -30
rect 169 -38 172 -32
rect 178 -38 183 -32
rect 169 -40 183 -38
rect 117 -46 127 -44
rect 82 -49 92 -47
rect 49 -56 72 -51
rect 49 -58 55 -56
rect 66 -58 72 -56
rect 82 -54 84 -49
rect 90 -54 92 -49
rect 82 -56 92 -54
rect 101 -48 111 -46
rect 101 -54 103 -48
rect 109 -54 111 -48
rect 138 -51 144 -40
rect 101 -56 111 -54
rect 82 -58 88 -56
rect 105 -58 111 -56
rect 121 -56 144 -51
rect 121 -58 127 -56
rect 138 -58 144 -56
rect 177 -58 183 -40
rect 194 -43 200 -29
rect 240 -30 246 -24
rect 232 -32 246 -30
rect 232 -38 235 -32
rect 241 -38 246 -32
rect 232 -40 246 -38
rect 194 -45 208 -43
rect 194 -51 200 -45
rect 206 -51 208 -45
rect 194 -53 208 -51
rect 240 -49 246 -40
rect 257 -43 263 -24
rect 302 -30 308 -24
rect 294 -32 308 -30
rect 294 -38 297 -32
rect 303 -38 308 -32
rect 294 -40 308 -38
rect 257 -45 271 -43
rect 257 -49 263 -45
rect 194 -58 200 -53
rect 240 -54 249 -49
rect 243 -58 249 -54
rect 254 -51 263 -49
rect 269 -51 271 -45
rect 254 -53 271 -51
rect 302 -49 308 -40
rect 319 -43 325 -24
rect 319 -45 333 -43
rect 319 -49 325 -45
rect 254 -55 263 -53
rect 302 -54 311 -49
rect 254 -58 260 -55
rect 305 -58 311 -54
rect 316 -51 325 -49
rect 331 -51 333 -45
rect 316 -53 333 -51
rect 316 -55 325 -53
rect 316 -58 322 -55
rect 49 -97 55 -92
rect 66 -97 72 -92
rect 82 -97 88 -92
rect 105 -97 111 -92
rect 121 -97 127 -92
rect 138 -97 144 -92
rect 177 -97 183 -92
rect 194 -97 200 -92
rect 243 -97 249 -92
rect 254 -97 260 -92
rect 305 -97 311 -92
rect 316 -97 322 -92
<< polycontact >>
rect 33 62 39 68
rect 55 62 61 68
rect 72 62 78 68
rect 27 46 33 52
rect 62 46 68 52
rect 93 46 99 52
rect 142 46 148 52
rect 170 59 176 65
rect 205 46 211 52
rect 233 59 239 65
rect 307 63 313 68
rect 326 62 332 68
rect 277 46 283 52
rect 302 42 308 48
rect 342 53 348 58
rect 357 46 363 52
rect 54 -38 60 -32
rect 79 -34 85 -28
rect 119 -44 125 -39
rect 134 -38 140 -32
rect 172 -38 178 -32
rect 84 -54 90 -49
rect 103 -54 109 -48
rect 235 -38 241 -32
rect 200 -51 206 -45
rect 297 -38 303 -32
rect 263 -51 269 -45
rect 325 -51 331 -45
<< metal1 >>
rect 0 120 387 127
rect 0 115 11 120
rect 16 115 35 120
rect 40 115 59 120
rect 64 115 83 120
rect 88 115 107 120
rect 112 115 139 120
rect 144 115 163 120
rect 168 115 202 120
rect 207 115 226 120
rect 231 115 264 120
rect 269 115 288 120
rect 293 115 312 120
rect 317 115 336 120
rect 341 115 360 120
rect 365 115 387 120
rect 0 113 387 115
rect 11 104 16 106
rect 11 68 16 96
rect 28 104 33 113
rect 61 104 66 106
rect 28 94 33 96
rect 60 96 61 97
rect 60 91 66 96
rect 94 104 99 113
rect 94 94 99 96
rect 111 104 116 106
rect 60 83 66 85
rect 111 78 116 96
rect 55 73 116 78
rect 55 68 61 73
rect 11 62 33 68
rect 39 62 48 68
rect 11 36 16 62
rect 42 52 48 62
rect 70 62 72 68
rect 78 62 80 68
rect 55 60 61 62
rect 25 46 27 52
rect 33 46 35 52
rect 42 46 62 52
rect 68 46 70 52
rect 91 46 93 52
rect 99 46 101 52
rect 60 39 66 41
rect 11 21 16 23
rect 28 36 33 38
rect 60 30 61 33
rect 28 14 33 23
rect 61 21 66 23
rect 94 36 99 38
rect 94 14 99 23
rect 111 36 116 73
rect 142 104 147 113
rect 170 104 175 106
rect 170 79 175 81
rect 156 78 175 79
rect 142 72 147 74
rect 154 72 156 78
rect 162 74 175 78
rect 202 104 207 113
rect 219 104 224 106
rect 219 78 224 79
rect 236 104 241 113
rect 162 72 164 74
rect 202 72 207 74
rect 217 72 219 78
rect 225 72 227 78
rect 236 72 241 74
rect 264 104 269 106
rect 281 104 286 113
rect 317 104 322 106
rect 317 93 322 99
rect 316 91 322 93
rect 353 104 358 113
rect 314 85 316 91
rect 322 85 324 91
rect 281 78 286 80
rect 140 46 142 52
rect 148 46 150 52
rect 111 21 116 23
rect 139 36 144 38
rect 139 14 144 23
rect 156 36 161 72
rect 168 59 170 65
rect 176 59 178 65
rect 203 46 205 52
rect 211 46 213 52
rect 156 21 161 23
rect 173 36 178 38
rect 219 37 224 72
rect 264 67 269 74
rect 307 75 347 80
rect 353 78 358 80
rect 370 104 375 106
rect 307 68 313 75
rect 342 70 347 75
rect 370 70 375 74
rect 326 68 332 70
rect 231 59 233 65
rect 239 59 241 65
rect 264 62 300 67
rect 305 63 307 68
rect 313 63 315 68
rect 173 14 178 23
rect 205 32 224 37
rect 233 36 238 38
rect 205 29 210 32
rect 205 21 210 23
rect 233 14 238 23
rect 264 36 269 62
rect 294 58 300 62
rect 326 58 332 62
rect 342 64 375 70
rect 342 59 348 64
rect 294 53 332 58
rect 340 58 350 59
rect 340 53 342 58
rect 348 53 350 58
rect 275 46 277 52
rect 283 46 285 52
rect 355 48 357 52
rect 300 42 302 48
rect 308 46 357 48
rect 363 46 365 52
rect 308 42 362 46
rect 264 21 269 23
rect 281 36 286 38
rect 316 36 322 37
rect 314 30 316 36
rect 322 30 324 36
rect 353 35 358 37
rect 316 28 322 30
rect 281 14 286 23
rect 317 21 322 23
rect 353 14 358 23
rect 370 36 375 64
rect 370 21 375 23
rect 0 12 387 14
rect 0 2 11 12
rect 16 2 35 12
rect 40 2 59 12
rect 64 2 83 12
rect 88 2 107 12
rect 112 2 139 12
rect 144 2 163 12
rect 168 2 202 12
rect 207 2 226 12
rect 231 2 264 12
rect 269 2 288 12
rect 293 7 312 12
rect 317 7 336 12
rect 341 7 360 12
rect 365 7 387 12
rect 293 2 387 7
rect 0 0 387 2
rect 41 -9 46 -7
rect 41 -48 46 -22
rect 58 -9 63 0
rect 94 -9 99 -7
rect 93 -16 99 -14
rect 130 -9 135 0
rect 91 -22 93 -16
rect 99 -22 101 -16
rect 58 -24 63 -22
rect 93 -23 99 -22
rect 130 -23 135 -21
rect 147 -9 152 -7
rect 52 -38 54 -32
rect 60 -38 62 -32
rect 77 -34 79 -28
rect 85 -32 139 -28
rect 85 -34 134 -32
rect 132 -38 134 -34
rect 140 -38 142 -32
rect 71 -44 109 -39
rect 71 -48 77 -44
rect 41 -53 77 -48
rect 103 -48 109 -44
rect 117 -44 119 -39
rect 125 -44 127 -39
rect 117 -45 127 -44
rect 41 -60 46 -53
rect 82 -54 84 -49
rect 90 -54 92 -49
rect 84 -61 90 -54
rect 103 -56 109 -54
rect 119 -50 125 -45
rect 147 -50 152 -22
rect 172 -9 177 -7
rect 172 -18 177 -15
rect 200 -9 205 0
rect 172 -23 191 -18
rect 170 -38 172 -32
rect 178 -38 180 -32
rect 119 -56 152 -50
rect 119 -61 124 -56
rect 41 -92 46 -90
rect 58 -66 63 -64
rect 84 -66 124 -61
rect 147 -60 152 -56
rect 186 -58 191 -23
rect 200 -24 205 -22
rect 232 -9 237 0
rect 232 -24 237 -22
rect 249 -9 254 -7
rect 233 -38 235 -32
rect 241 -38 243 -32
rect 198 -51 200 -45
rect 206 -51 208 -45
rect 249 -58 254 -22
rect 266 -9 271 0
rect 266 -24 271 -22
rect 294 -9 299 0
rect 294 -24 299 -22
rect 311 -9 316 -7
rect 295 -38 297 -32
rect 303 -38 305 -32
rect 261 -51 263 -45
rect 269 -51 271 -45
rect 311 -58 316 -22
rect 328 -9 333 0
rect 328 -24 333 -22
rect 323 -51 325 -45
rect 331 -51 333 -45
rect 130 -66 135 -64
rect 91 -77 93 -71
rect 99 -77 101 -71
rect 93 -79 99 -77
rect 58 -99 63 -90
rect 94 -85 99 -79
rect 94 -92 99 -90
rect 130 -99 135 -90
rect 147 -92 152 -90
rect 169 -60 174 -58
rect 184 -64 186 -58
rect 192 -64 194 -58
rect 203 -60 208 -58
rect 169 -99 174 -90
rect 186 -65 191 -64
rect 186 -92 191 -90
rect 203 -99 208 -90
rect 235 -60 240 -58
rect 247 -64 249 -58
rect 255 -60 257 -58
rect 297 -60 302 -58
rect 255 -64 268 -60
rect 249 -65 268 -64
rect 235 -99 240 -90
rect 263 -67 268 -65
rect 263 -92 268 -90
rect 309 -64 311 -58
rect 317 -60 319 -58
rect 317 -64 330 -60
rect 311 -65 330 -64
rect 297 -99 302 -90
rect 325 -67 330 -65
rect 325 -92 330 -90
rect 0 -101 387 -99
rect 0 -106 41 -101
rect 46 -106 65 -101
rect 70 -106 89 -101
rect 94 -106 113 -101
rect 118 -106 137 -101
rect 142 -106 169 -101
rect 174 -106 193 -101
rect 198 -106 232 -101
rect 237 -106 256 -101
rect 261 -106 294 -101
rect 299 -106 318 -101
rect 323 -106 387 -101
rect 0 -113 387 -106
<< via1 >>
rect 60 85 66 91
rect 72 62 78 68
rect 27 46 33 52
rect 93 46 99 52
rect 60 37 66 39
rect 60 33 61 37
rect 61 33 66 37
rect 156 72 162 78
rect 219 72 225 78
rect 316 85 322 91
rect 142 46 148 52
rect 170 59 176 65
rect 205 46 211 52
rect 233 59 239 65
rect 277 46 283 52
rect 357 46 363 52
rect 316 30 322 36
rect 93 -22 99 -16
rect 54 -38 60 -32
rect 79 -34 85 -28
rect 134 -38 140 -32
rect 172 -38 178 -32
rect 235 -38 241 -32
rect 200 -51 206 -45
rect 297 -38 303 -32
rect 263 -51 269 -45
rect 325 -51 331 -45
rect 93 -77 99 -71
rect 186 -64 192 -58
rect 249 -64 255 -58
rect 311 -64 317 -58
<< metal2 >>
rect 60 92 66 97
rect 316 92 322 93
rect 59 91 67 92
rect 315 91 323 92
rect 59 85 60 91
rect 66 85 148 91
rect 59 84 67 85
rect 59 83 66 84
rect 27 53 33 54
rect 26 52 34 53
rect 26 46 27 52
rect 33 46 34 52
rect 26 45 34 46
rect 27 26 33 45
rect 59 40 65 83
rect 72 69 79 70
rect 71 68 80 69
rect 71 62 72 68
rect 78 62 113 68
rect 71 61 80 62
rect 72 60 80 61
rect 58 39 68 40
rect 58 33 60 39
rect 66 33 68 39
rect 58 32 68 33
rect 74 26 80 60
rect 93 53 99 54
rect 92 52 100 53
rect 107 52 113 62
rect 142 65 148 85
rect 315 85 316 91
rect 322 85 323 91
rect 315 84 323 85
rect 154 78 164 79
rect 154 72 156 78
rect 162 72 164 78
rect 154 71 164 72
rect 217 78 227 79
rect 217 72 219 78
rect 225 72 227 78
rect 217 71 227 72
rect 168 65 178 66
rect 231 65 241 66
rect 142 59 170 65
rect 176 59 233 65
rect 239 59 241 65
rect 168 58 178 59
rect 231 58 241 59
rect 140 52 150 53
rect 91 46 93 52
rect 99 46 101 52
rect 107 46 142 52
rect 148 46 150 52
rect 92 45 100 46
rect 140 45 150 46
rect 203 52 213 53
rect 276 52 284 53
rect 203 46 205 52
rect 211 46 213 52
rect 275 46 277 52
rect 283 46 285 52
rect 203 45 213 46
rect 276 45 284 46
rect 27 20 80 26
rect 27 -2 33 20
rect 93 9 99 45
rect 316 37 322 84
rect 356 52 364 53
rect 355 46 357 52
rect 363 46 365 52
rect 356 45 364 46
rect 314 36 324 37
rect 314 30 316 36
rect 322 30 324 36
rect 314 29 324 30
rect 8 -8 33 -2
rect 39 3 99 9
rect 39 -14 45 3
rect 8 -20 45 -14
rect 54 -9 178 -3
rect 54 -31 60 -9
rect 91 -16 101 -15
rect 91 -22 93 -16
rect 99 -22 101 -16
rect 91 -23 101 -22
rect 78 -28 86 -27
rect 53 -32 61 -31
rect 8 -38 54 -32
rect 60 -38 62 -32
rect 78 -34 79 -28
rect 85 -34 86 -28
rect 78 -35 86 -34
rect 53 -39 61 -38
rect 79 -45 85 -35
rect 8 -51 85 -45
rect 93 -45 99 -23
rect 172 -31 178 -9
rect 133 -32 141 -31
rect 170 -32 180 -31
rect 132 -38 134 -32
rect 140 -38 142 -32
rect 170 -38 172 -32
rect 178 -38 180 -32
rect 133 -39 141 -38
rect 170 -39 180 -38
rect 233 -32 243 -31
rect 233 -38 235 -32
rect 241 -38 243 -32
rect 233 -39 243 -38
rect 295 -32 305 -31
rect 295 -38 297 -32
rect 303 -38 305 -32
rect 295 -39 305 -38
rect 198 -45 208 -44
rect 93 -51 200 -45
rect 206 -51 208 -45
rect 93 -70 99 -51
rect 198 -52 208 -51
rect 261 -45 271 -44
rect 261 -51 263 -45
rect 269 -51 271 -45
rect 261 -52 271 -51
rect 323 -45 333 -44
rect 323 -51 325 -45
rect 331 -51 333 -45
rect 323 -52 333 -51
rect 184 -58 194 -57
rect 184 -64 186 -58
rect 192 -64 194 -58
rect 184 -65 194 -64
rect 247 -58 257 -57
rect 247 -64 249 -58
rect 255 -64 257 -58
rect 247 -65 257 -64
rect 309 -58 319 -57
rect 309 -64 311 -58
rect 317 -64 319 -58
rect 309 -65 319 -64
rect 92 -71 100 -70
rect 92 -77 93 -71
rect 99 -77 100 -71
rect 92 -78 100 -77
rect 93 -79 99 -78
<< labels >>
rlabel metal1 13 117 13 117 1 my_nxor_0.VDD
rlabel psubdiffcont 13 9 13 9 1 my_nxor_0.VSS
rlabel psubdiffcont 13 4 13 4 5 my_xor_0.VSS
rlabel psubdiffcont 141 5 141 5 5 my_nand_0.VSS
rlabel psubdiffcont 141 9 141 9 1 my_nor_0.VSS
rlabel nsubdiffcont 141 117 141 117 1 my_nor_0.VDD
rlabel via1 159 75 159 75 1 my_nor_0.Y
rlabel via1 173 62 173 62 1 my_nor_0.B
rlabel via1 145 49 145 49 1 my_nor_0.A
rlabel psubdiffcont 204 5 204 5 5 my_nor_0.VSS
rlabel psubdiffcont 204 9 204 9 1 my_nand_0.VSS
rlabel nsubdiffcont 204 118 204 118 1 my_nand_0.VDD
rlabel psubdiffcont 266 5 266 5 5 my_nor_0.VSS
rlabel via1 280 49 280 49 1 my_xor_0.A
rlabel via1 360 49 360 49 1 my_xor_0.B
rlabel via1 319 87 319 87 1 my_xor_0.Y
rlabel nsubdiffcont 266 118 266 118 1 my_xor_0.VDD
rlabel psubdiffcont 266 10 266 10 1 my_xor_0.VSS
rlabel metal2 30 49 30 49 1 my_nxor_0.A
rlabel via1 57 -35 57 -35 5 my_xor_0.A
rlabel via1 137 -35 137 -35 5 my_xor_0.B
rlabel via1 96 -73 96 -73 5 my_xor_0.Y
rlabel nsubdiffcont 43 -104 43 -104 5 my_xor_0.VDD
rlabel via1 175 -35 175 -35 5 my_nand_0.A
rlabel via1 203 -48 203 -48 5 my_nand_0.B
rlabel via1 189 -61 189 -61 5 my_nand_0.Y
rlabel nsubdiffcont 171 -104 171 -104 5 my_nand_0.VDD
rlabel via1 238 -35 238 -35 5 my_nor_0.A
rlabel via1 266 -48 266 -48 5 my_nor_0.B
rlabel via1 252 -61 252 -61 5 my_nor_0.Y
rlabel nsubdiffcont 234 -103 234 -103 5 my_nor_0.VDD
rlabel nsubdiffcont 296 -103 296 -103 5 my_nor_0.VDD
rlabel via1 314 -61 314 -61 5 my_nor_0.Y
rlabel via1 328 -48 328 -48 5 my_nor_0.B
rlabel via1 300 -35 300 -35 5 my_nor_0.A
rlabel metal2 63 87 63 87 1 my_nxor_0.Y
rlabel metal2 96 49 96 49 1 my_nxor_0.B
rlabel via1 222 75 222 75 1 my_nand_0.Y
rlabel via1 236 62 236 62 1 my_nand_0_A
rlabel via1 208 49 208 49 1 my_nand_0_B
<< end >>
