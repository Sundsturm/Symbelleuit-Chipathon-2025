VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 2bit_comp_1x
  CLASS BLOCK ;
  FOREIGN 2bit_comp_1x ;
  ORIGIN 0.000 5.650 ;
  SIZE 19.600 BY 12.000 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 0.000 -4.950 19.600 -2.450 ;
        RECT 0.900 -5.650 18.650 -4.950 ;
      LAYER Metal1 ;
        RECT 2.300 -4.950 2.550 -3.200 ;
        RECT 5.900 -4.950 6.150 -3.200 ;
        RECT 8.250 -4.950 8.500 -2.900 ;
        RECT 9.950 -4.950 10.200 -2.900 ;
        RECT 11.600 -4.950 11.850 -2.900 ;
        RECT 15.550 -4.950 15.800 -2.900 ;
        RECT 0.000 -5.650 19.600 -4.950 ;
    END
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 19.600 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 19.600 6.350 ;
        RECT 1.400 4.700 1.650 5.650 ;
        RECT 4.700 4.700 4.950 5.650 ;
        RECT 7.200 3.600 7.450 5.650 ;
        RECT 10.250 3.600 10.500 5.650 ;
        RECT 11.950 3.600 12.200 5.650 ;
        RECT 14.300 3.900 14.550 5.650 ;
        RECT 17.900 3.900 18.150 5.650 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.700 0.700 4.950 1.900 ;
        RECT 7.050 0.700 7.300 1.900 ;
        RECT 8.750 0.700 9.000 1.900 ;
        RECT 11.800 0.700 12.050 1.900 ;
        RECT 14.300 0.700 14.550 1.900 ;
        RECT 17.900 0.700 18.150 1.850 ;
        RECT 0.000 0.000 19.600 0.700 ;
        RECT 2.300 -1.200 2.550 0.000 ;
        RECT 5.900 -1.150 6.150 0.000 ;
        RECT 9.800 -1.200 10.050 0.000 ;
        RECT 11.450 -1.200 11.700 0.000 ;
        RECT 13.150 -1.200 13.400 0.000 ;
        RECT 15.400 -1.200 15.650 0.000 ;
        RECT 17.100 -1.200 17.350 0.000 ;
    END
  END VSS
  PIN B0
    USE SIGNAL ;
    ANTENNAGATEAREA 2.550000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 -1.900 2.500 -1.600 ;
        RECT 8.300 -1.900 8.800 -1.600 ;
      LAYER Metal2 ;
        RECT 2.100 -0.450 7.100 -0.150 ;
        RECT 2.100 -1.550 2.400 -0.450 ;
        RECT 6.800 -1.300 7.100 -0.450 ;
        RECT 6.800 -1.550 8.700 -1.300 ;
        RECT 2.050 -1.600 2.450 -1.550 ;
        RECT 6.800 -1.600 8.800 -1.550 ;
        RECT 2.000 -1.900 2.500 -1.600 ;
        RECT 2.050 -1.950 2.450 -1.900 ;
        RECT 8.300 -1.950 8.800 -1.600 ;
    END
  END B0
  PIN A0
    USE SIGNAL ;
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 -1.600 6.350 -1.400 ;
        RECT 3.250 -1.700 6.500 -1.600 ;
        RECT 6.000 -1.900 6.500 -1.700 ;
      LAYER Metal2 ;
        RECT 6.050 -1.600 6.450 -1.550 ;
        RECT 6.000 -1.900 6.500 -1.600 ;
        RECT 6.050 -1.950 6.450 -1.900 ;
    END
  END A0
  PIN B1
    USE SIGNAL ;
    ANTENNAGATEAREA 2.805000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 3.100 4.000 3.400 ;
        RECT 8.500 2.950 9.000 3.250 ;
        RECT 1.250 2.300 1.750 2.600 ;
      LAYER Metal2 ;
        RECT 3.600 3.450 3.950 3.500 ;
        RECT 3.550 3.400 4.000 3.450 ;
        RECT 3.550 3.250 7.500 3.400 ;
        RECT 8.500 3.250 9.000 3.300 ;
        RECT 3.550 3.100 9.000 3.250 ;
        RECT 3.550 3.050 4.000 3.100 ;
        RECT 3.600 3.000 4.000 3.050 ;
        RECT 1.350 2.650 1.650 2.700 ;
        RECT 1.300 2.250 1.700 2.650 ;
        RECT 1.350 1.300 1.650 2.250 ;
        RECT 3.700 1.300 4.000 3.000 ;
        RECT 7.200 2.950 9.000 3.100 ;
        RECT 8.500 2.900 9.000 2.950 ;
        RECT 1.350 1.000 4.000 1.300 ;
    END
  END B1
  PIN A1
    USE SIGNAL ;
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 2.300 5.050 2.600 ;
      LAYER Metal2 ;
        RECT 4.650 2.650 4.950 2.700 ;
        RECT 4.600 2.600 5.000 2.650 ;
        RECT 4.550 2.300 5.050 2.600 ;
        RECT 4.600 2.250 5.000 2.300 ;
        RECT 4.650 2.200 4.950 2.250 ;
    END
  END A1
  PIN L
    USE SIGNAL ;
    ANTENNAGATEAREA 1.275000 ;
    ANTENNADIFFAREA 2.167500 ;
    PORT
      LAYER Metal1 ;
        RECT 16.100 4.650 16.350 5.300 ;
        RECT 16.050 4.550 16.350 4.650 ;
        RECT 15.950 4.250 16.450 4.550 ;
        RECT 16.050 1.800 16.350 1.850 ;
        RECT 15.950 1.500 16.450 1.800 ;
        RECT 16.050 1.400 16.350 1.500 ;
        RECT 16.100 1.050 16.350 1.400 ;
        RECT 15.450 -1.900 15.950 -1.600 ;
      LAYER Metal2 ;
        RECT 16.050 4.600 16.350 4.650 ;
        RECT 16.000 4.550 16.400 4.600 ;
        RECT 16.000 4.250 19.150 4.550 ;
        RECT 16.000 4.200 16.400 4.250 ;
        RECT 16.050 1.850 16.350 4.200 ;
        RECT 15.950 1.450 16.450 1.850 ;
        RECT 15.450 -1.600 15.950 -1.550 ;
        RECT 18.800 -1.600 19.150 4.250 ;
        RECT 15.450 -1.900 19.150 -1.600 ;
        RECT 15.450 -1.950 15.950 -1.900 ;
    END
  END L
  PIN G
    USE SIGNAL ;
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal1 ;
        RECT 16.250 -2.900 16.500 -0.350 ;
        RECT 16.150 -3.000 16.650 -2.900 ;
        RECT 16.150 -3.200 17.200 -3.000 ;
        RECT 16.250 -3.250 17.200 -3.200 ;
        RECT 16.950 -4.600 17.200 -3.250 ;
      LAYER Metal2 ;
        RECT 16.150 -3.250 16.650 -2.850 ;
    END
  END G
  PIN E
    USE SIGNAL ;
    ANTENNAGATEAREA 1.275000 ;
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal1 ;
        RECT 12.300 -2.900 12.550 -0.350 ;
        RECT 16.850 -2.550 17.350 -2.250 ;
        RECT 12.200 -3.000 12.700 -2.900 ;
        RECT 12.200 -3.200 13.250 -3.000 ;
        RECT 12.300 -3.250 13.250 -3.200 ;
        RECT 13.000 -4.600 13.250 -3.250 ;
      LAYER Metal2 ;
        RECT 16.850 -2.250 17.350 -2.200 ;
        RECT 14.650 -2.550 17.350 -2.250 ;
        RECT 12.200 -2.900 12.700 -2.850 ;
        RECT 14.650 -2.900 14.950 -2.550 ;
        RECT 16.850 -2.600 17.350 -2.550 ;
        RECT 12.200 -3.200 14.950 -2.900 ;
        RECT 12.200 -3.250 12.700 -3.200 ;
    END
  END E
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.400 0.800 5.300 ;
        RECT 3.050 4.850 3.300 5.300 ;
        RECT 3.000 4.150 3.300 4.850 ;
        RECT 5.550 3.900 5.800 5.300 ;
        RECT 6.250 4.750 6.650 5.250 ;
        RECT 6.200 4.000 6.600 4.500 ;
        RECT 2.750 3.650 5.800 3.900 ;
        RECT 0.550 3.100 2.400 3.400 ;
        RECT 0.550 1.050 0.800 3.100 ;
        RECT 2.100 2.600 2.400 3.100 ;
        RECT 2.750 3.000 3.050 3.650 ;
        RECT 2.100 2.300 3.500 2.600 ;
        RECT 3.000 1.500 3.300 2.050 ;
        RECT 3.050 1.050 3.300 1.500 ;
        RECT 5.550 1.050 5.800 3.650 ;
        RECT 6.250 2.600 6.550 4.000 ;
        RECT 8.600 3.950 8.850 5.300 ;
        RECT 9.400 4.750 9.800 5.250 ;
        RECT 7.900 3.900 8.850 3.950 ;
        RECT 11.100 3.900 11.350 5.300 ;
        RECT 7.800 3.700 8.850 3.900 ;
        RECT 7.800 3.600 8.300 3.700 ;
        RECT 11.000 3.600 11.500 3.900 ;
        RECT 6.250 2.300 7.600 2.600 ;
        RECT 7.900 1.050 8.150 3.600 ;
        RECT 10.300 2.300 10.800 2.600 ;
        RECT 11.100 1.850 11.350 3.600 ;
        RECT 13.450 3.350 13.700 5.300 ;
        RECT 15.600 3.750 17.600 4.000 ;
        RECT 15.600 3.400 15.900 3.750 ;
        RECT 17.350 3.500 17.600 3.750 ;
        RECT 18.750 3.500 19.000 5.300 ;
        RECT 11.700 2.950 12.200 3.250 ;
        RECT 13.450 3.100 15.250 3.350 ;
        RECT 15.500 3.150 16.000 3.400 ;
        RECT 9.450 1.200 9.850 1.700 ;
        RECT 10.400 1.600 11.350 1.850 ;
        RECT 10.400 1.050 10.650 1.600 ;
        RECT 12.600 1.200 13.000 1.700 ;
        RECT 13.450 1.050 13.700 3.100 ;
        RECT 14.950 2.900 15.250 3.100 ;
        RECT 16.550 2.900 16.850 3.500 ;
        RECT 17.350 3.200 19.000 3.500 ;
        RECT 17.350 2.950 17.650 3.200 ;
        RECT 14.950 2.650 16.850 2.900 ;
        RECT 17.250 2.650 17.750 2.950 ;
        RECT 14.000 2.300 14.500 2.600 ;
        RECT 18.000 2.400 18.500 2.600 ;
        RECT 15.250 2.300 18.500 2.400 ;
        RECT 15.250 2.100 18.350 2.300 ;
        RECT 18.750 1.050 19.000 3.200 ;
        RECT 1.450 -2.400 1.700 -0.350 ;
        RECT 4.100 -0.700 4.350 -0.350 ;
        RECT 4.050 -0.800 4.350 -0.700 ;
        RECT 3.950 -1.100 4.450 -0.800 ;
        RECT 4.050 -1.150 4.350 -1.100 ;
        RECT 2.950 -2.200 4.850 -1.950 ;
        RECT 2.950 -2.400 3.250 -2.200 ;
        RECT 1.450 -2.650 3.250 -2.400 ;
        RECT 1.450 -4.600 1.700 -2.650 ;
        RECT 3.500 -2.700 4.000 -2.450 ;
        RECT 3.600 -3.050 3.900 -2.700 ;
        RECT 4.550 -2.800 4.850 -2.200 ;
        RECT 5.250 -2.250 5.750 -1.950 ;
        RECT 5.350 -2.500 5.650 -2.250 ;
        RECT 6.750 -2.500 7.000 -0.350 ;
        RECT 7.450 -1.000 7.850 -0.500 ;
        RECT 8.400 -0.900 8.650 -0.350 ;
        RECT 8.400 -1.150 9.350 -0.900 ;
        RECT 10.600 -1.000 11.000 -0.500 ;
        RECT 5.350 -2.800 7.000 -2.500 ;
        RECT 5.350 -3.050 5.600 -2.800 ;
        RECT 3.600 -3.300 5.600 -3.050 ;
        RECT 3.950 -3.850 4.450 -3.550 ;
        RECT 4.050 -3.950 4.350 -3.850 ;
        RECT 4.100 -4.600 4.350 -3.950 ;
        RECT 6.750 -4.600 7.000 -2.800 ;
        RECT 9.100 -2.900 9.350 -1.150 ;
        RECT 11.500 -1.900 12.000 -1.600 ;
        RECT 9.700 -2.550 10.200 -2.250 ;
        RECT 12.900 -2.550 13.400 -2.250 ;
        RECT 9.000 -3.200 9.500 -2.900 ;
        RECT 9.100 -4.600 9.350 -3.200 ;
        RECT 10.650 -4.550 11.050 -4.050 ;
        RECT 13.800 -4.550 14.200 -4.050 ;
        RECT 14.600 -4.550 15.000 -4.050 ;
        RECT 17.750 -4.550 18.150 -4.050 ;
      LAYER Metal2 ;
        RECT 3.000 4.600 3.300 4.850 ;
        RECT 6.200 4.800 9.850 5.200 ;
        RECT 10.400 4.850 14.400 5.150 ;
        RECT 2.950 4.500 3.350 4.600 ;
        RECT 10.400 4.500 10.700 4.850 ;
        RECT 2.950 4.200 6.600 4.500 ;
        RECT 2.950 4.150 3.300 4.200 ;
        RECT 2.950 2.000 3.250 4.150 ;
        RECT 6.200 4.000 6.600 4.200 ;
        RECT 7.900 4.200 10.700 4.500 ;
        RECT 7.900 3.950 8.300 4.200 ;
        RECT 7.800 3.550 8.300 3.950 ;
        RECT 11.000 3.550 11.500 3.950 ;
        RECT 11.700 3.250 12.200 3.300 ;
        RECT 11.700 2.950 13.700 3.250 ;
        RECT 11.700 2.900 12.200 2.950 ;
        RECT 7.100 2.600 7.600 2.650 ;
        RECT 10.300 2.600 10.800 2.650 ;
        RECT 7.100 2.300 10.800 2.600 ;
        RECT 7.100 2.250 7.600 2.300 ;
        RECT 10.300 2.250 10.800 2.300 ;
        RECT 2.900 1.600 3.400 2.000 ;
        RECT 9.400 1.600 9.900 1.650 ;
        RECT 12.550 1.600 13.050 1.650 ;
        RECT 9.400 1.300 13.050 1.600 ;
        RECT 9.400 1.250 9.900 1.300 ;
        RECT 12.550 1.250 13.050 1.300 ;
        RECT 13.400 1.150 13.700 2.950 ;
        RECT 14.100 2.650 14.400 4.850 ;
        RECT 14.050 2.600 14.450 2.650 ;
        RECT 18.050 2.600 18.450 2.650 ;
        RECT 14.000 2.300 14.500 2.600 ;
        RECT 18.000 2.300 18.500 2.600 ;
        RECT 14.050 2.250 14.450 2.300 ;
        RECT 18.050 2.250 18.450 2.300 ;
        RECT 18.100 1.150 18.400 2.250 ;
        RECT 13.400 0.850 18.400 1.150 ;
        RECT 7.400 -0.600 7.900 -0.550 ;
        RECT 10.550 -0.600 11.050 -0.550 ;
        RECT 3.950 -1.150 4.450 -0.750 ;
        RECT 7.400 -0.900 11.050 -0.600 ;
        RECT 7.400 -0.950 7.900 -0.900 ;
        RECT 10.550 -0.950 11.050 -0.900 ;
        RECT 4.050 -3.500 4.350 -1.150 ;
        RECT 11.500 -1.600 12.000 -1.550 ;
        RECT 13.400 -1.600 13.700 0.850 ;
        RECT 11.500 -1.900 13.700 -1.600 ;
        RECT 11.500 -1.950 12.000 -1.900 ;
        RECT 9.700 -2.250 10.200 -2.200 ;
        RECT 12.900 -2.250 13.400 -2.200 ;
        RECT 7.600 -2.550 13.400 -2.250 ;
        RECT 4.000 -3.550 4.400 -3.500 ;
        RECT 7.600 -3.550 7.900 -2.550 ;
        RECT 9.700 -2.600 10.200 -2.550 ;
        RECT 12.900 -2.600 13.400 -2.550 ;
        RECT 9.000 -3.250 9.500 -2.850 ;
        RECT 4.000 -3.850 7.900 -3.550 ;
        RECT 4.000 -3.900 4.400 -3.850 ;
        RECT 4.050 -3.950 4.350 -3.900 ;
        RECT 10.600 -4.500 14.250 -4.100 ;
        RECT 14.550 -4.500 18.200 -4.100 ;
      LAYER Metal3 ;
        RECT 11.700 3.250 12.200 3.350 ;
        RECT 9.100 2.950 12.200 3.250 ;
        RECT 9.100 -2.800 9.400 2.950 ;
        RECT 11.700 2.850 12.200 2.950 ;
        RECT 9.000 -3.300 9.500 -2.800 ;
  END
END 2bit_comp_1x
END LIBRARY

