magic
tech gf180mcuD
magscale 1 5
timestamp 1755595404
<< error_p >>
rect 820 420 858 423
<< nwell >>
rect 0 315 1960 635
rect 0 -495 1960 -245
rect 90 -565 1865 -495
<< nmos >>
rect 95 105 125 190
rect 180 105 210 190
rect 245 105 275 190
rect 360 105 390 190
rect 425 105 455 190
rect 510 105 540 190
rect 745 105 775 190
rect 830 105 860 190
rect 995 105 1025 190
rect 1080 105 1110 190
rect 1135 105 1165 190
rect 1220 105 1250 190
rect 1385 105 1415 190
rect 1470 105 1500 190
rect 1550 105 1580 190
rect 1665 105 1695 190
rect 1745 105 1775 190
rect 1830 105 1860 190
rect 185 -120 215 -35
rect 270 -120 300 -35
rect 350 -120 380 -35
rect 465 -120 495 -35
rect 545 -120 575 -35
rect 630 -120 660 -35
rect 795 -120 825 -35
rect 880 -120 910 -35
rect 935 -120 965 -35
rect 1020 -120 1050 -35
rect 1185 -120 1215 -35
rect 1270 -120 1300 -35
rect 1580 -120 1610 -35
rect 1665 -120 1695 -35
<< pmos >>
rect 95 360 125 530
rect 180 360 210 530
rect 245 360 275 530
rect 360 360 390 530
rect 425 360 455 530
rect 510 360 540 530
rect 675 360 705 530
rect 760 360 790 530
rect 815 360 845 530
rect 900 360 930 530
rect 1065 360 1095 530
rect 1150 360 1180 530
rect 1385 360 1415 530
rect 1470 360 1500 530
rect 1550 360 1580 530
rect 1665 360 1695 530
rect 1745 360 1775 530
rect 1830 360 1860 530
rect 185 -460 215 -290
rect 270 -460 300 -290
rect 350 -460 380 -290
rect 465 -460 495 -290
rect 545 -460 575 -290
rect 630 -460 660 -290
rect 865 -460 895 -290
rect 950 -460 980 -290
rect 1115 -460 1145 -290
rect 1200 -460 1230 -290
rect 1255 -460 1285 -290
rect 1340 -460 1370 -290
rect 1510 -460 1540 -290
rect 1595 -460 1625 -290
rect 1650 -460 1680 -290
rect 1735 -460 1765 -290
<< ndiff >>
rect 290 190 340 195
rect 45 180 95 190
rect 45 115 55 180
rect 80 115 95 180
rect 45 105 95 115
rect 125 180 180 190
rect 125 115 140 180
rect 165 115 180 180
rect 125 105 180 115
rect 210 105 245 190
rect 275 185 360 190
rect 275 115 305 185
rect 330 115 360 185
rect 275 105 360 115
rect 390 105 425 190
rect 455 180 510 190
rect 455 115 470 180
rect 495 115 510 180
rect 455 105 510 115
rect 540 180 590 190
rect 540 115 555 180
rect 580 115 590 180
rect 540 105 590 115
rect 695 180 745 190
rect 695 115 705 180
rect 730 115 745 180
rect 695 105 745 115
rect 775 180 830 190
rect 775 115 790 180
rect 815 115 830 180
rect 775 105 830 115
rect 860 180 910 190
rect 860 115 875 180
rect 900 115 910 180
rect 860 105 910 115
rect 940 160 995 190
rect 940 130 950 160
rect 980 130 995 160
rect 940 105 995 130
rect 1025 145 1080 190
rect 1025 115 1040 145
rect 1065 115 1080 145
rect 1025 105 1080 115
rect 1110 105 1135 190
rect 1165 180 1220 190
rect 1165 115 1180 180
rect 1205 115 1220 180
rect 1165 105 1220 115
rect 1250 160 1305 190
rect 1250 130 1265 160
rect 1295 130 1305 160
rect 1250 105 1305 130
rect 1335 180 1385 190
rect 1335 115 1345 180
rect 1370 115 1385 180
rect 1335 105 1385 115
rect 1415 180 1470 190
rect 1415 115 1430 180
rect 1455 115 1470 180
rect 1415 105 1470 115
rect 1500 105 1550 190
rect 1580 140 1665 190
rect 1580 115 1610 140
rect 1635 115 1665 140
rect 1580 105 1665 115
rect 1695 105 1745 190
rect 1775 175 1830 190
rect 1775 115 1790 175
rect 1815 115 1830 175
rect 1775 105 1830 115
rect 1860 180 1910 190
rect 1860 115 1875 180
rect 1900 115 1910 180
rect 1860 105 1910 115
rect 135 -45 185 -35
rect 135 -110 145 -45
rect 170 -110 185 -45
rect 135 -120 185 -110
rect 215 -45 270 -35
rect 215 -110 230 -45
rect 255 -110 270 -45
rect 215 -120 270 -110
rect 300 -120 350 -35
rect 380 -45 465 -35
rect 380 -70 410 -45
rect 435 -70 465 -45
rect 380 -120 465 -70
rect 495 -120 545 -35
rect 575 -45 630 -35
rect 575 -105 590 -45
rect 615 -105 630 -45
rect 575 -120 630 -105
rect 660 -45 710 -35
rect 660 -110 675 -45
rect 700 -110 710 -45
rect 660 -120 710 -110
rect 740 -60 795 -35
rect 740 -90 750 -60
rect 780 -90 795 -60
rect 740 -120 795 -90
rect 825 -45 880 -35
rect 825 -75 840 -45
rect 865 -75 880 -45
rect 825 -120 880 -75
rect 910 -120 935 -35
rect 965 -45 1020 -35
rect 965 -110 980 -45
rect 1005 -110 1020 -45
rect 965 -120 1020 -110
rect 1050 -60 1105 -35
rect 1050 -90 1065 -60
rect 1095 -90 1105 -60
rect 1050 -120 1105 -90
rect 1135 -45 1185 -35
rect 1135 -110 1145 -45
rect 1170 -110 1185 -45
rect 1135 -120 1185 -110
rect 1215 -45 1270 -35
rect 1215 -110 1230 -45
rect 1255 -110 1270 -45
rect 1215 -120 1270 -110
rect 1300 -45 1350 -35
rect 1300 -110 1315 -45
rect 1340 -110 1350 -45
rect 1300 -120 1350 -110
rect 1530 -45 1580 -35
rect 1530 -110 1540 -45
rect 1565 -110 1580 -45
rect 1530 -120 1580 -110
rect 1610 -45 1665 -35
rect 1610 -110 1625 -45
rect 1650 -110 1665 -45
rect 1610 -120 1665 -110
rect 1695 -45 1745 -35
rect 1695 -110 1710 -45
rect 1735 -110 1745 -45
rect 1695 -120 1745 -110
<< pdiff >>
rect 45 520 95 530
rect 45 480 55 520
rect 80 480 95 520
rect 45 360 95 480
rect 125 520 180 530
rect 125 480 140 520
rect 165 480 180 520
rect 125 360 180 480
rect 210 360 245 530
rect 275 520 360 530
rect 275 480 305 520
rect 330 480 360 520
rect 275 360 360 480
rect 390 360 425 530
rect 455 520 510 530
rect 455 480 470 520
rect 495 480 510 520
rect 455 360 510 480
rect 540 520 590 530
rect 540 480 555 520
rect 580 480 590 520
rect 540 360 590 480
rect 620 515 675 530
rect 620 485 630 515
rect 660 485 675 515
rect 620 360 675 485
rect 705 520 760 530
rect 705 370 720 520
rect 745 370 760 520
rect 705 360 760 370
rect 790 360 815 530
rect 845 520 900 530
rect 845 405 860 520
rect 885 405 900 520
rect 845 360 900 405
rect 930 515 985 530
rect 930 485 945 515
rect 975 485 985 515
rect 930 360 985 485
rect 1015 520 1065 530
rect 1015 370 1025 520
rect 1050 370 1065 520
rect 1015 360 1065 370
rect 1095 520 1150 530
rect 1095 395 1110 520
rect 1135 395 1150 520
rect 1095 360 1150 395
rect 1180 520 1230 530
rect 1180 370 1195 520
rect 1220 370 1230 520
rect 1180 360 1230 370
rect 1335 520 1385 530
rect 1335 370 1345 520
rect 1370 370 1385 520
rect 1335 360 1385 370
rect 1415 520 1470 530
rect 1415 400 1430 520
rect 1455 400 1470 520
rect 1415 360 1470 400
rect 1500 360 1550 530
rect 1580 520 1665 530
rect 1580 495 1610 520
rect 1635 495 1665 520
rect 1580 360 1665 495
rect 1695 360 1745 530
rect 1775 520 1830 530
rect 1775 400 1790 520
rect 1815 400 1830 520
rect 1775 360 1830 400
rect 1860 520 1910 530
rect 1860 370 1875 520
rect 1900 370 1910 520
rect 1860 360 1910 370
rect 135 -300 185 -290
rect 135 -450 145 -300
rect 170 -450 185 -300
rect 135 -460 185 -450
rect 215 -330 270 -290
rect 215 -450 230 -330
rect 255 -450 270 -330
rect 215 -460 270 -450
rect 300 -460 350 -290
rect 380 -425 465 -290
rect 380 -450 410 -425
rect 435 -450 465 -425
rect 380 -460 465 -450
rect 495 -460 545 -290
rect 575 -330 630 -290
rect 575 -450 590 -330
rect 615 -450 630 -330
rect 575 -460 630 -450
rect 660 -300 710 -290
rect 660 -450 675 -300
rect 700 -450 710 -300
rect 660 -460 710 -450
rect 815 -300 865 -290
rect 815 -450 825 -300
rect 850 -450 865 -300
rect 815 -460 865 -450
rect 895 -325 950 -290
rect 895 -450 910 -325
rect 935 -450 950 -325
rect 895 -460 950 -450
rect 980 -300 1030 -290
rect 980 -450 995 -300
rect 1020 -450 1030 -300
rect 980 -460 1030 -450
rect 1060 -415 1115 -290
rect 1060 -445 1070 -415
rect 1100 -445 1115 -415
rect 1060 -460 1115 -445
rect 1145 -300 1200 -290
rect 1145 -450 1160 -300
rect 1185 -450 1200 -300
rect 1145 -460 1200 -450
rect 1230 -460 1255 -290
rect 1285 -335 1340 -290
rect 1285 -450 1300 -335
rect 1325 -450 1340 -335
rect 1285 -460 1340 -450
rect 1370 -415 1425 -290
rect 1370 -445 1385 -415
rect 1415 -445 1425 -415
rect 1370 -460 1425 -445
rect 1455 -415 1510 -290
rect 1455 -445 1465 -415
rect 1495 -445 1510 -415
rect 1455 -460 1510 -445
rect 1540 -300 1595 -290
rect 1540 -450 1555 -300
rect 1580 -450 1595 -300
rect 1540 -460 1595 -450
rect 1625 -460 1650 -290
rect 1680 -335 1735 -290
rect 1680 -450 1695 -335
rect 1720 -450 1735 -335
rect 1680 -460 1735 -450
rect 1765 -415 1820 -290
rect 1765 -445 1780 -415
rect 1810 -445 1820 -415
rect 1765 -460 1820 -445
<< ndiffc >>
rect 55 115 80 180
rect 140 115 165 180
rect 305 115 330 185
rect 470 115 495 180
rect 555 115 580 180
rect 705 115 730 180
rect 790 115 815 180
rect 875 115 900 180
rect 950 130 980 160
rect 1040 115 1065 145
rect 1180 115 1205 180
rect 1265 130 1295 160
rect 1345 115 1370 180
rect 1430 115 1455 180
rect 1610 115 1635 140
rect 1790 115 1815 175
rect 1875 115 1900 180
rect 145 -110 170 -45
rect 230 -110 255 -45
rect 410 -70 435 -45
rect 590 -105 615 -45
rect 675 -110 700 -45
rect 750 -90 780 -60
rect 840 -75 865 -45
rect 980 -110 1005 -45
rect 1065 -90 1095 -60
rect 1145 -110 1170 -45
rect 1230 -110 1255 -45
rect 1315 -110 1340 -45
rect 1540 -110 1565 -45
rect 1625 -110 1650 -45
rect 1710 -110 1735 -45
<< pdiffc >>
rect 55 480 80 520
rect 140 480 165 520
rect 305 480 330 520
rect 470 480 495 520
rect 555 480 580 520
rect 630 485 660 515
rect 720 370 745 520
rect 860 405 885 520
rect 945 485 975 515
rect 1025 370 1050 520
rect 1110 395 1135 520
rect 1195 370 1220 520
rect 1345 370 1370 520
rect 1430 400 1455 520
rect 1610 495 1635 520
rect 1790 400 1815 520
rect 1875 370 1900 520
rect 145 -450 170 -300
rect 230 -450 255 -330
rect 410 -450 435 -425
rect 590 -450 615 -330
rect 675 -450 700 -300
rect 825 -450 850 -300
rect 910 -450 935 -325
rect 995 -450 1020 -300
rect 1070 -445 1100 -415
rect 1160 -450 1185 -300
rect 1300 -450 1325 -335
rect 1385 -445 1415 -415
rect 1465 -445 1495 -415
rect 1555 -450 1580 -300
rect 1695 -450 1720 -335
rect 1780 -445 1810 -415
<< psubdiff >>
rect 115 50 190 60
rect 115 20 140 50
rect 165 20 190 50
rect 115 10 190 20
rect 285 50 360 60
rect 285 20 310 50
rect 335 20 360 50
rect 285 10 360 20
rect 445 50 520 60
rect 445 20 470 50
rect 495 20 520 50
rect 445 10 520 20
rect 565 50 640 60
rect 565 20 590 50
rect 615 20 640 50
rect 565 10 640 20
rect 680 50 755 60
rect 680 20 705 50
rect 730 20 755 50
rect 680 10 755 20
rect 850 50 925 60
rect 850 20 875 50
rect 900 20 925 50
rect 850 10 925 20
rect 955 50 1030 60
rect 955 20 980 50
rect 1005 20 1030 50
rect 955 10 1030 20
rect 1140 50 1215 60
rect 1140 20 1165 50
rect 1190 20 1215 50
rect 1140 10 1215 20
rect 1290 50 1365 60
rect 1290 20 1315 50
rect 1340 20 1365 50
rect 1290 10 1365 20
rect 1515 50 1590 60
rect 1515 20 1540 50
rect 1565 20 1590 50
rect 1515 10 1590 20
rect 1685 50 1760 60
rect 1685 20 1710 50
rect 1735 20 1760 50
rect 1685 10 1760 20
rect 1835 50 1910 60
rect 1835 20 1860 50
rect 1885 20 1910 50
rect 1835 10 1910 20
<< nsubdiff >>
rect 30 600 105 610
rect 30 575 55 600
rect 80 575 105 600
rect 30 565 105 575
rect 150 600 225 610
rect 150 575 175 600
rect 200 575 225 600
rect 150 565 225 575
rect 270 600 345 610
rect 270 575 295 600
rect 320 575 345 600
rect 270 565 345 575
rect 390 600 465 610
rect 390 575 415 600
rect 440 575 465 600
rect 390 565 465 575
rect 510 600 585 610
rect 510 575 535 600
rect 560 575 585 600
rect 510 565 585 575
rect 680 600 755 610
rect 680 575 705 600
rect 730 575 755 600
rect 680 565 755 575
rect 800 600 875 610
rect 800 575 825 600
rect 850 575 875 600
rect 800 565 875 575
rect 1000 600 1075 610
rect 1000 575 1025 600
rect 1050 575 1075 600
rect 1000 565 1075 575
rect 1120 600 1195 610
rect 1120 575 1145 600
rect 1170 575 1195 600
rect 1120 565 1195 575
rect 1320 600 1395 610
rect 1320 575 1345 600
rect 1370 575 1395 600
rect 1320 565 1395 575
rect 1440 600 1515 610
rect 1440 575 1465 600
rect 1490 575 1515 600
rect 1440 565 1515 575
rect 1560 600 1635 610
rect 1560 575 1585 600
rect 1610 575 1635 600
rect 1560 565 1635 575
rect 1680 600 1755 610
rect 1680 575 1705 600
rect 1730 575 1755 600
rect 1680 565 1755 575
rect 1800 600 1875 610
rect 1800 575 1825 600
rect 1850 575 1875 600
rect 1800 565 1875 575
rect 120 -505 195 -495
rect 120 -530 145 -505
rect 170 -530 195 -505
rect 120 -540 195 -530
rect 240 -505 315 -495
rect 240 -530 265 -505
rect 290 -530 315 -505
rect 240 -540 315 -530
rect 360 -505 435 -495
rect 360 -530 385 -505
rect 410 -530 435 -505
rect 360 -540 435 -530
rect 480 -505 555 -495
rect 480 -530 505 -505
rect 530 -530 555 -505
rect 480 -540 555 -530
rect 600 -505 675 -495
rect 600 -530 625 -505
rect 650 -530 675 -505
rect 600 -540 675 -530
rect 800 -505 875 -495
rect 800 -530 825 -505
rect 850 -530 875 -505
rect 800 -540 875 -530
rect 920 -505 995 -495
rect 920 -530 945 -505
rect 970 -530 995 -505
rect 920 -540 995 -530
rect 1120 -505 1195 -495
rect 1120 -530 1145 -505
rect 1170 -530 1195 -505
rect 1120 -540 1195 -530
rect 1240 -505 1315 -495
rect 1240 -530 1265 -505
rect 1290 -530 1315 -505
rect 1240 -540 1315 -530
rect 1515 -505 1590 -495
rect 1515 -530 1540 -505
rect 1565 -530 1590 -505
rect 1515 -540 1590 -530
rect 1635 -505 1710 -495
rect 1635 -530 1660 -505
rect 1685 -530 1710 -505
rect 1635 -540 1710 -530
<< psubdiffcont >>
rect 140 20 165 50
rect 310 20 335 50
rect 470 20 495 50
rect 590 20 615 50
rect 705 20 730 50
rect 875 20 900 50
rect 980 20 1005 50
rect 1165 20 1190 50
rect 1315 20 1340 50
rect 1540 20 1565 50
rect 1710 20 1735 50
rect 1860 20 1885 50
<< nsubdiffcont >>
rect 55 575 80 600
rect 175 575 200 600
rect 295 575 320 600
rect 415 575 440 600
rect 535 575 560 600
rect 705 575 730 600
rect 825 575 850 600
rect 1025 575 1050 600
rect 1145 575 1170 600
rect 1345 575 1370 600
rect 1465 575 1490 600
rect 1585 575 1610 600
rect 1705 575 1730 600
rect 1825 575 1850 600
rect 145 -530 170 -505
rect 265 -530 290 -505
rect 385 -530 410 -505
rect 505 -530 530 -505
rect 625 -530 650 -505
rect 825 -530 850 -505
rect 945 -530 970 -505
rect 1145 -530 1170 -505
rect 1265 -530 1290 -505
rect 1540 -530 1565 -505
rect 1660 -530 1685 -505
<< polysilicon >>
rect 95 530 125 555
rect 180 530 210 555
rect 245 530 275 555
rect 360 530 390 555
rect 425 530 455 555
rect 510 530 540 555
rect 675 530 705 555
rect 760 530 790 555
rect 815 530 845 555
rect 900 530 930 555
rect 1065 530 1095 555
rect 1150 530 1180 555
rect 1385 530 1415 555
rect 1470 530 1500 555
rect 1550 530 1580 555
rect 1665 530 1695 555
rect 1745 530 1775 555
rect 1830 530 1860 555
rect 95 270 125 360
rect 180 350 210 360
rect 155 340 210 350
rect 155 310 165 340
rect 195 310 210 340
rect 155 300 210 310
rect 245 350 275 360
rect 360 350 390 360
rect 425 350 455 360
rect 510 350 540 360
rect 245 340 315 350
rect 245 310 275 340
rect 305 310 315 340
rect 245 300 315 310
rect 350 340 400 350
rect 350 310 360 340
rect 390 310 400 340
rect 425 325 540 350
rect 350 300 400 310
rect 95 260 175 270
rect 95 230 135 260
rect 165 255 175 260
rect 165 230 210 255
rect 95 220 210 230
rect 95 190 125 220
rect 180 190 210 220
rect 245 190 275 300
rect 510 270 540 325
rect 675 340 705 360
rect 760 340 790 360
rect 675 315 790 340
rect 815 345 845 360
rect 815 335 860 345
rect 900 335 930 360
rect 815 325 930 335
rect 815 315 860 325
rect 745 270 775 315
rect 300 260 350 270
rect 455 260 540 270
rect 300 230 310 260
rect 340 230 390 260
rect 455 245 465 260
rect 300 220 390 230
rect 360 190 390 220
rect 425 230 465 245
rect 495 230 540 260
rect 425 220 540 230
rect 705 260 775 270
rect 705 230 720 260
rect 750 230 775 260
rect 705 220 775 230
rect 425 190 455 220
rect 510 190 540 220
rect 745 190 775 220
rect 830 295 860 315
rect 890 305 930 325
rect 890 295 900 305
rect 830 285 900 295
rect 830 190 860 285
rect 1065 270 1095 360
rect 1020 260 1095 270
rect 1020 230 1040 260
rect 1070 230 1095 260
rect 1020 220 1095 230
rect 995 200 1040 220
rect 1065 215 1095 220
rect 1150 335 1180 360
rect 1385 350 1415 360
rect 1470 350 1500 360
rect 1150 325 1220 335
rect 1150 295 1180 325
rect 1210 295 1220 325
rect 1150 285 1220 295
rect 1385 325 1500 350
rect 1550 350 1580 360
rect 1665 350 1695 360
rect 1550 340 1600 350
rect 1150 225 1180 285
rect 1385 270 1415 325
rect 1550 315 1560 340
rect 1590 315 1600 340
rect 1550 305 1600 315
rect 1645 340 1695 350
rect 1645 310 1655 340
rect 1685 310 1695 340
rect 1745 350 1775 360
rect 1830 350 1860 360
rect 1745 325 1860 350
rect 1645 300 1695 310
rect 1385 260 1450 270
rect 1385 230 1410 260
rect 1440 230 1450 260
rect 1150 215 1250 225
rect 1065 200 1110 215
rect 995 190 1025 200
rect 1080 190 1110 200
rect 1135 200 1250 215
rect 1135 190 1165 200
rect 1220 190 1250 200
rect 1385 220 1450 230
rect 1525 240 1580 250
rect 1385 200 1500 220
rect 1525 210 1535 240
rect 1565 210 1580 240
rect 1525 200 1580 210
rect 1385 190 1415 200
rect 1470 190 1500 200
rect 1550 190 1580 200
rect 1665 190 1695 300
rect 1725 290 1775 300
rect 1725 265 1735 290
rect 1765 265 1775 290
rect 1830 270 1860 325
rect 1725 255 1775 265
rect 1745 190 1775 255
rect 1800 260 1860 270
rect 1800 230 1810 260
rect 1840 230 1860 260
rect 1800 220 1860 230
rect 1830 190 1860 220
rect 95 80 125 105
rect 180 80 210 105
rect 245 80 275 105
rect 360 80 390 105
rect 425 80 455 105
rect 510 80 540 105
rect 745 80 775 105
rect 830 80 860 105
rect 995 80 1025 105
rect 1080 80 1110 105
rect 1135 80 1165 105
rect 1220 80 1250 105
rect 1385 80 1415 105
rect 1470 80 1500 105
rect 1550 80 1580 105
rect 1665 80 1695 105
rect 1745 80 1775 105
rect 1830 80 1860 105
rect 185 -35 215 -10
rect 270 -35 300 -10
rect 350 -35 380 -10
rect 465 -35 495 -10
rect 545 -35 575 -10
rect 630 -35 660 -10
rect 795 -35 825 -10
rect 880 -35 910 -10
rect 935 -35 965 -10
rect 1020 -35 1050 -10
rect 1185 -35 1215 -10
rect 1270 -35 1300 -10
rect 1580 -35 1610 -10
rect 1665 -35 1695 -10
rect 185 -130 215 -120
rect 270 -130 300 -120
rect 350 -130 380 -120
rect 185 -150 300 -130
rect 325 -140 380 -130
rect 185 -160 250 -150
rect 185 -190 210 -160
rect 240 -190 250 -160
rect 325 -170 335 -140
rect 365 -170 380 -140
rect 325 -180 380 -170
rect 185 -200 250 -190
rect 185 -255 215 -200
rect 465 -230 495 -120
rect 545 -185 575 -120
rect 630 -150 660 -120
rect 795 -130 825 -120
rect 880 -130 910 -120
rect 795 -150 840 -130
rect 865 -145 910 -130
rect 935 -130 965 -120
rect 1020 -130 1050 -120
rect 935 -145 1050 -130
rect 865 -150 895 -145
rect 525 -195 575 -185
rect 525 -220 535 -195
rect 565 -220 575 -195
rect 600 -160 660 -150
rect 600 -190 610 -160
rect 640 -190 660 -160
rect 600 -200 660 -190
rect 820 -160 895 -150
rect 820 -190 840 -160
rect 870 -190 895 -160
rect 820 -200 895 -190
rect 525 -230 575 -220
rect 350 -245 400 -235
rect 185 -280 300 -255
rect 185 -290 215 -280
rect 270 -290 300 -280
rect 350 -270 360 -245
rect 390 -270 400 -245
rect 350 -280 400 -270
rect 445 -240 495 -230
rect 445 -270 455 -240
rect 485 -270 495 -240
rect 630 -255 660 -200
rect 445 -280 495 -270
rect 350 -290 380 -280
rect 465 -290 495 -280
rect 545 -280 660 -255
rect 545 -290 575 -280
rect 630 -290 660 -280
rect 865 -290 895 -200
rect 950 -155 1050 -145
rect 1185 -150 1215 -120
rect 950 -215 980 -155
rect 1145 -160 1215 -150
rect 1145 -190 1160 -160
rect 1190 -190 1215 -160
rect 1145 -200 1215 -190
rect 950 -225 1020 -215
rect 950 -255 980 -225
rect 1010 -255 1020 -225
rect 1185 -245 1215 -200
rect 1270 -215 1300 -120
rect 1580 -150 1610 -120
rect 1540 -160 1610 -150
rect 1540 -190 1555 -160
rect 1585 -190 1610 -160
rect 1540 -200 1610 -190
rect 1270 -225 1340 -215
rect 1270 -245 1300 -225
rect 950 -265 1020 -255
rect 950 -290 980 -265
rect 1115 -270 1230 -245
rect 1115 -290 1145 -270
rect 1200 -290 1230 -270
rect 1255 -255 1300 -245
rect 1330 -235 1340 -225
rect 1330 -255 1370 -235
rect 1580 -245 1610 -200
rect 1665 -215 1695 -120
rect 1665 -225 1735 -215
rect 1665 -245 1695 -225
rect 1255 -265 1370 -255
rect 1255 -275 1300 -265
rect 1255 -290 1285 -275
rect 1340 -290 1370 -265
rect 1510 -270 1625 -245
rect 1510 -290 1540 -270
rect 1595 -290 1625 -270
rect 1650 -255 1695 -245
rect 1725 -235 1735 -225
rect 1725 -255 1765 -235
rect 1650 -265 1765 -255
rect 1650 -275 1695 -265
rect 1650 -290 1680 -275
rect 1735 -290 1765 -265
rect 185 -485 215 -460
rect 270 -485 300 -460
rect 350 -485 380 -460
rect 465 -485 495 -460
rect 545 -485 575 -460
rect 630 -485 660 -460
rect 865 -485 895 -460
rect 950 -485 980 -460
rect 1115 -485 1145 -460
rect 1200 -485 1230 -460
rect 1255 -485 1285 -460
rect 1340 -485 1370 -460
rect 1510 -485 1540 -460
rect 1595 -485 1625 -460
rect 1650 -485 1680 -460
rect 1735 -485 1765 -460
<< polycontact >>
rect 165 310 195 340
rect 275 310 305 340
rect 360 310 390 340
rect 135 230 165 260
rect 310 230 340 260
rect 465 230 495 260
rect 720 230 750 260
rect 860 295 890 325
rect 1040 230 1070 260
rect 1180 295 1210 325
rect 1560 315 1590 340
rect 1655 310 1685 340
rect 1410 230 1440 260
rect 1535 210 1565 240
rect 1735 265 1765 290
rect 1810 230 1840 260
rect 210 -190 240 -160
rect 335 -170 365 -140
rect 535 -220 565 -195
rect 610 -190 640 -160
rect 840 -190 870 -160
rect 360 -270 390 -245
rect 455 -270 485 -240
rect 1160 -190 1190 -160
rect 980 -255 1010 -225
rect 1555 -190 1585 -160
rect 1300 -255 1330 -225
rect 1695 -255 1725 -225
<< metal1 >>
rect 0 600 1960 635
rect 0 575 55 600
rect 80 575 175 600
rect 200 575 295 600
rect 320 575 415 600
rect 440 575 535 600
rect 560 575 705 600
rect 730 575 825 600
rect 850 575 1025 600
rect 1050 575 1145 600
rect 1170 575 1345 600
rect 1370 575 1465 600
rect 1490 575 1585 600
rect 1610 575 1705 600
rect 1730 575 1825 600
rect 1850 575 1960 600
rect 0 565 1960 575
rect 55 520 80 530
rect 55 340 80 480
rect 140 520 165 565
rect 305 520 330 530
rect 140 470 165 480
rect 300 480 305 485
rect 300 455 330 480
rect 470 520 495 565
rect 470 470 495 480
rect 555 520 580 530
rect 300 415 330 425
rect 555 390 580 480
rect 625 515 665 525
rect 625 485 630 515
rect 660 485 665 515
rect 625 475 665 485
rect 720 520 745 565
rect 620 440 660 450
rect 620 410 625 440
rect 655 410 660 440
rect 620 400 660 410
rect 275 365 580 390
rect 275 340 305 365
rect 55 310 165 340
rect 195 310 240 340
rect 55 180 80 310
rect 210 260 240 310
rect 350 310 360 340
rect 390 310 400 340
rect 275 300 305 310
rect 125 230 135 260
rect 165 230 175 260
rect 210 230 310 260
rect 340 230 350 260
rect 455 230 465 260
rect 495 230 505 260
rect 300 195 330 205
rect 55 105 80 115
rect 140 180 165 190
rect 300 150 305 165
rect 140 70 165 115
rect 305 105 330 115
rect 470 180 495 190
rect 470 70 495 115
rect 555 180 580 365
rect 625 260 655 400
rect 860 520 885 530
rect 940 515 980 525
rect 940 485 945 515
rect 975 485 980 515
rect 940 475 980 485
rect 1025 520 1050 565
rect 860 395 885 405
rect 790 390 885 395
rect 720 360 745 370
rect 780 360 790 390
rect 820 370 885 390
rect 1110 520 1135 530
rect 1110 390 1135 395
rect 1195 520 1220 565
rect 820 360 830 370
rect 1025 360 1050 370
rect 1100 360 1110 390
rect 1140 360 1150 390
rect 1195 360 1220 370
rect 1345 520 1370 530
rect 1430 520 1455 565
rect 1610 520 1635 530
rect 1610 465 1635 495
rect 1605 455 1635 465
rect 1790 520 1815 565
rect 1595 425 1605 455
rect 1635 425 1645 455
rect 1430 390 1455 400
rect 625 230 720 260
rect 750 230 760 260
rect 555 105 580 115
rect 705 180 730 190
rect 705 70 730 115
rect 790 180 815 360
rect 850 295 860 325
rect 890 295 900 325
rect 1030 230 1040 260
rect 1070 230 1080 260
rect 790 105 815 115
rect 875 180 900 190
rect 1110 185 1135 360
rect 1345 335 1370 370
rect 1560 375 1760 400
rect 1790 390 1815 400
rect 1875 520 1900 530
rect 1560 340 1590 375
rect 1735 350 1760 375
rect 1875 350 1900 370
rect 1655 340 1685 350
rect 1170 295 1180 325
rect 1210 295 1220 325
rect 1345 310 1525 335
rect 1550 315 1560 340
rect 1590 315 1600 340
rect 945 160 985 170
rect 945 130 950 160
rect 980 130 985 160
rect 945 120 985 130
rect 1040 160 1135 185
rect 1180 180 1205 190
rect 1040 145 1065 160
rect 875 70 900 115
rect 1040 105 1065 115
rect 1345 180 1370 310
rect 1495 290 1525 310
rect 1655 290 1685 310
rect 1735 320 1900 350
rect 1735 295 1765 320
rect 1495 265 1685 290
rect 1725 290 1775 295
rect 1725 265 1735 290
rect 1765 265 1775 290
rect 1400 230 1410 260
rect 1440 230 1450 260
rect 1800 240 1810 260
rect 1525 210 1535 240
rect 1565 230 1810 240
rect 1840 230 1850 260
rect 1565 210 1835 230
rect 1260 160 1300 170
rect 1260 130 1265 160
rect 1295 130 1300 160
rect 1260 120 1300 130
rect 1180 70 1205 115
rect 1345 105 1370 115
rect 1430 180 1455 190
rect 1605 180 1635 185
rect 1595 150 1605 180
rect 1635 150 1645 180
rect 1790 175 1815 185
rect 1605 140 1635 150
rect 1430 70 1455 115
rect 1610 105 1635 115
rect 1790 70 1815 115
rect 1875 180 1900 320
rect 1875 105 1900 115
rect 0 50 1960 70
rect 0 20 140 50
rect 165 20 310 50
rect 335 20 470 50
rect 495 20 590 50
rect 615 20 705 50
rect 730 20 875 50
rect 900 20 980 50
rect 1005 20 1165 50
rect 1190 20 1315 50
rect 1340 20 1540 50
rect 1565 20 1710 50
rect 1735 20 1860 50
rect 1885 20 1960 50
rect 0 0 1960 20
rect 145 -45 170 -35
rect 145 -240 170 -110
rect 230 -45 255 0
rect 410 -45 435 -35
rect 405 -80 435 -70
rect 590 -45 615 0
rect 395 -110 405 -80
rect 435 -110 445 -80
rect 230 -120 255 -110
rect 405 -115 435 -110
rect 590 -115 615 -105
rect 675 -45 700 -35
rect 840 -45 865 -35
rect 745 -60 785 -50
rect 745 -90 750 -60
rect 780 -90 785 -60
rect 745 -100 785 -90
rect 840 -90 865 -75
rect 980 -45 1005 0
rect 200 -190 210 -160
rect 240 -190 250 -160
rect 325 -170 335 -140
rect 365 -160 635 -140
rect 365 -170 610 -160
rect 600 -190 610 -170
rect 640 -190 650 -160
rect 295 -220 485 -195
rect 295 -240 325 -220
rect 145 -265 325 -240
rect 455 -240 485 -220
rect 525 -220 535 -195
rect 565 -220 575 -195
rect 525 -225 575 -220
rect 145 -300 170 -265
rect 350 -270 360 -245
rect 390 -270 400 -245
rect 360 -305 390 -270
rect 455 -280 485 -270
rect 535 -250 565 -225
rect 675 -250 700 -110
rect 840 -115 935 -90
rect 830 -190 840 -160
rect 870 -190 880 -160
rect 535 -280 700 -250
rect 535 -305 560 -280
rect 145 -460 170 -450
rect 230 -330 255 -320
rect 360 -330 560 -305
rect 675 -300 700 -280
rect 910 -290 935 -115
rect 1145 -45 1170 0
rect 1060 -60 1100 -50
rect 1060 -90 1065 -60
rect 1095 -90 1100 -60
rect 1060 -100 1100 -90
rect 980 -120 1005 -110
rect 1145 -120 1170 -110
rect 1230 -45 1255 -35
rect 1150 -190 1160 -160
rect 1190 -190 1200 -160
rect 970 -255 980 -225
rect 1010 -255 1020 -225
rect 1230 -290 1255 -110
rect 1315 -45 1340 0
rect 1315 -120 1340 -110
rect 1540 -45 1565 0
rect 1540 -120 1565 -110
rect 1625 -45 1650 -35
rect 1545 -190 1555 -160
rect 1585 -190 1595 -160
rect 1290 -255 1300 -225
rect 1330 -255 1340 -225
rect 1625 -290 1650 -110
rect 1710 -45 1735 0
rect 1710 -120 1735 -110
rect 1685 -255 1695 -225
rect 1725 -255 1735 -225
rect 590 -330 615 -320
rect 395 -385 405 -355
rect 435 -385 445 -355
rect 405 -395 435 -385
rect 230 -495 255 -450
rect 410 -425 435 -395
rect 410 -460 435 -450
rect 590 -495 615 -450
rect 675 -460 700 -450
rect 825 -300 850 -290
rect 900 -320 910 -290
rect 940 -320 950 -290
rect 995 -300 1020 -290
rect 825 -495 850 -450
rect 910 -325 935 -320
rect 910 -460 935 -450
rect 1160 -300 1185 -290
rect 995 -495 1020 -450
rect 1065 -415 1105 -405
rect 1065 -445 1070 -415
rect 1100 -445 1105 -415
rect 1065 -455 1105 -445
rect 1220 -320 1230 -290
rect 1260 -300 1270 -290
rect 1555 -300 1580 -290
rect 1260 -320 1325 -300
rect 1230 -325 1325 -320
rect 1160 -495 1185 -450
rect 1300 -335 1325 -325
rect 1300 -460 1325 -450
rect 1380 -415 1420 -405
rect 1380 -445 1385 -415
rect 1415 -445 1420 -415
rect 1380 -455 1420 -445
rect 1460 -415 1500 -405
rect 1460 -445 1465 -415
rect 1495 -445 1500 -415
rect 1460 -455 1500 -445
rect 1615 -320 1625 -290
rect 1655 -300 1665 -290
rect 1655 -320 1720 -300
rect 1625 -325 1720 -320
rect 1555 -495 1580 -450
rect 1695 -335 1720 -325
rect 1695 -460 1720 -450
rect 1775 -415 1815 -405
rect 1775 -445 1780 -415
rect 1810 -445 1815 -415
rect 1775 -455 1815 -445
rect 0 -505 1960 -495
rect 0 -530 145 -505
rect 170 -530 265 -505
rect 290 -530 385 -505
rect 410 -530 505 -505
rect 530 -530 625 -505
rect 650 -530 825 -505
rect 850 -530 945 -505
rect 970 -530 1145 -505
rect 1170 -530 1265 -505
rect 1290 -530 1540 -505
rect 1565 -530 1660 -505
rect 1685 -530 1960 -505
rect 0 -565 1960 -530
<< via1 >>
rect 300 425 330 455
rect 630 485 660 515
rect 625 410 655 440
rect 360 310 390 340
rect 135 230 165 260
rect 465 230 495 260
rect 300 185 330 195
rect 300 165 305 185
rect 305 165 330 185
rect 945 485 975 515
rect 790 360 820 390
rect 1110 360 1140 390
rect 1605 425 1635 455
rect 720 230 750 260
rect 860 295 890 325
rect 1040 230 1070 260
rect 1180 295 1210 325
rect 950 130 980 160
rect 1410 230 1440 260
rect 1810 230 1840 260
rect 1265 130 1295 160
rect 1605 150 1635 180
rect 405 -110 435 -80
rect 750 -90 780 -60
rect 210 -190 240 -160
rect 610 -190 640 -160
rect 840 -190 870 -160
rect 1065 -90 1095 -60
rect 1160 -190 1190 -160
rect 980 -255 1010 -225
rect 1555 -190 1585 -160
rect 1300 -255 1330 -225
rect 1695 -255 1725 -225
rect 405 -385 435 -355
rect 910 -320 940 -290
rect 1070 -445 1100 -415
rect 1230 -320 1260 -290
rect 1385 -445 1415 -415
rect 1465 -445 1495 -415
rect 1625 -320 1655 -290
rect 1780 -445 1810 -415
<< metal2 >>
rect 620 515 985 520
rect 620 485 630 515
rect 660 485 945 515
rect 975 485 985 515
rect 300 460 330 485
rect 620 480 985 485
rect 1040 485 1440 515
rect 295 455 335 460
rect 295 425 300 455
rect 330 450 335 455
rect 1040 450 1070 485
rect 330 440 660 450
rect 330 425 625 440
rect 295 420 625 425
rect 295 415 330 420
rect 135 265 165 270
rect 130 260 170 265
rect 130 230 135 260
rect 165 230 170 260
rect 130 225 170 230
rect 135 130 165 225
rect 295 200 325 415
rect 620 410 625 420
rect 655 410 660 440
rect 620 400 660 410
rect 790 420 1070 450
rect 790 395 820 420
rect 780 390 830 395
rect 780 360 790 390
rect 820 360 830 390
rect 780 355 830 360
rect 1100 390 1150 395
rect 1100 360 1110 390
rect 1140 360 1150 390
rect 1100 355 1150 360
rect 360 345 395 350
rect 355 340 400 345
rect 355 310 360 340
rect 390 325 750 340
rect 850 325 900 330
rect 390 310 860 325
rect 355 305 400 310
rect 360 300 400 305
rect 290 195 340 200
rect 290 165 300 195
rect 330 165 340 195
rect 290 160 340 165
rect 370 130 400 300
rect 720 295 860 310
rect 890 295 900 325
rect 850 290 900 295
rect 1170 290 1175 330
rect 1215 325 1220 330
rect 1215 295 1370 325
rect 1215 290 1220 295
rect 465 265 495 270
rect 460 260 500 265
rect 710 260 760 265
rect 1030 260 1080 265
rect 455 230 465 260
rect 495 230 505 260
rect 710 230 720 260
rect 750 230 1040 260
rect 1070 230 1080 260
rect 460 225 500 230
rect 710 225 760 230
rect 1030 225 1080 230
rect 465 220 495 225
rect 135 100 400 130
rect 940 160 990 165
rect 1255 160 1305 165
rect 940 130 950 160
rect 980 130 1265 160
rect 1295 130 1305 160
rect 940 125 990 130
rect 1255 125 1305 130
rect 1340 115 1370 295
rect 1410 265 1440 485
rect 1605 460 1635 465
rect 1600 455 1640 460
rect 1600 425 1605 455
rect 1635 425 1915 455
rect 1600 420 1640 425
rect 1405 260 1445 265
rect 1400 230 1410 260
rect 1440 230 1450 260
rect 1405 225 1445 230
rect 1605 185 1635 420
rect 1805 260 1845 265
rect 1800 230 1810 260
rect 1840 230 1850 260
rect 1805 225 1845 230
rect 1595 180 1645 185
rect 1595 150 1605 180
rect 1635 150 1645 180
rect 1595 145 1645 150
rect 1810 115 1840 225
rect 1340 85 1840 115
rect 210 -45 710 -15
rect 210 -155 240 -45
rect 395 -80 445 -75
rect 395 -110 405 -80
rect 435 -110 445 -80
rect 395 -115 445 -110
rect 205 -160 245 -155
rect 200 -190 210 -160
rect 240 -190 250 -160
rect 205 -195 245 -190
rect 405 -350 435 -115
rect 680 -130 710 -45
rect 740 -60 790 -55
rect 1055 -60 1105 -55
rect 740 -90 750 -60
rect 780 -90 1065 -60
rect 1095 -90 1105 -60
rect 740 -95 790 -90
rect 1055 -95 1105 -90
rect 680 -155 870 -130
rect 605 -160 645 -155
rect 680 -160 880 -155
rect 600 -190 610 -160
rect 640 -190 650 -160
rect 830 -190 840 -160
rect 870 -190 880 -160
rect 605 -195 645 -190
rect 830 -195 880 -190
rect 1150 -160 1200 -155
rect 1340 -160 1370 85
rect 1150 -190 1160 -160
rect 1190 -190 1370 -160
rect 1545 -160 1595 -155
rect 1880 -160 1915 425
rect 1545 -190 1555 -160
rect 1585 -190 1915 -160
rect 1150 -195 1200 -190
rect 1545 -195 1595 -190
rect 970 -225 1020 -220
rect 1290 -225 1340 -220
rect 1685 -225 1735 -220
rect 760 -255 980 -225
rect 1010 -255 1300 -225
rect 1330 -255 1340 -225
rect 400 -355 440 -350
rect 760 -355 790 -255
rect 970 -260 1020 -255
rect 1290 -260 1340 -255
rect 1465 -255 1695 -225
rect 1725 -255 1735 -225
rect 900 -325 905 -285
rect 945 -325 950 -285
rect 1220 -290 1270 -285
rect 1465 -290 1495 -255
rect 1685 -260 1735 -255
rect 1220 -320 1230 -290
rect 1260 -320 1495 -290
rect 1615 -290 1665 -285
rect 1615 -320 1625 -290
rect 1655 -320 1665 -290
rect 1220 -325 1270 -320
rect 1615 -325 1665 -320
rect 400 -385 405 -355
rect 435 -385 790 -355
rect 400 -390 440 -385
rect 405 -395 435 -390
rect 1060 -415 1425 -410
rect 1060 -445 1070 -415
rect 1100 -445 1385 -415
rect 1415 -445 1425 -415
rect 1060 -450 1425 -445
rect 1455 -415 1820 -410
rect 1455 -445 1465 -415
rect 1495 -445 1780 -415
rect 1810 -445 1820 -415
rect 1455 -450 1820 -445
<< via2 >>
rect 1175 325 1215 330
rect 1175 295 1180 325
rect 1180 295 1210 325
rect 1210 295 1215 325
rect 1175 290 1215 295
rect 905 -290 945 -285
rect 905 -320 910 -290
rect 910 -320 940 -290
rect 940 -320 945 -290
rect 905 -325 945 -320
<< metal3 >>
rect 1170 330 1220 335
rect 1170 325 1175 330
rect 910 295 1175 325
rect 910 -280 940 295
rect 1170 290 1175 295
rect 1215 290 1220 330
rect 1170 285 1220 290
rect 900 -285 950 -280
rect 900 -325 905 -285
rect 945 -325 950 -285
rect 900 -330 950 -325
<< labels >>
rlabel metal2 150 245 150 245 1 my_nxor_0.A
rlabel metal2 315 435 315 435 1 my_nxor_0.Y
rlabel metal2 480 245 480 245 1 my_nxor_0.B
rlabel via1 805 375 805 375 1 my_nor_0.Y
rlabel metal2 1055 245 1055 245 1 my_nand_0.A
rlabel via2 1195 310 1195 310 1 my_nand_0.B
rlabel metal2 1125 375 1125 375 1 my_nand_0.Y
rlabel via1 420 -365 420 -365 5 my_xor_0.Y
rlabel via1 625 -175 625 -175 5 my_xor_0.B
rlabel via1 225 -175 225 -175 5 my_xor_0.A
rlabel via1 1175 -175 1175 -175 1 my_nor_1.A
rlabel via1 1315 -240 1315 -240 1 my_nor_1.B
rlabel via1 1245 -305 1245 -305 1 my_nor_1.Y
rlabel via1 1570 -175 1570 -175 1 my_nor_2.A
rlabel via1 1710 -240 1710 -240 1 my_nor_2.B
rlabel via1 1640 -305 1640 -305 1 my_nor_2.Y
rlabel via1 1425 245 1425 245 1 my_xor_1.A
rlabel via1 1825 245 1825 245 1 my_xor_1.B
rlabel via1 1620 440 1620 440 1 my_xor_1.Y
rlabel via1 855 -175 855 -175 1 my_nand_1.A
rlabel via1 995 -240 995 -240 1 my_nand_1.B
rlabel via1 925 -305 925 -305 1 my_nand_1.Y
rlabel metal1 15 -530 15 -530 1 VDD
rlabel metal1 20 605 20 605 1 VDD
rlabel metal1 20 35 20 35 1 VSS
rlabel via1 150 235 150 235 1 B1
rlabel via1 480 235 480 235 1 A1
rlabel via1 225 -170 225 -170 1 B0
rlabel via1 625 -170 625 -170 1 A0
rlabel via1 735 245 735 245 1 my_nor_0.B
rlabel via1 875 310 875 310 1 my_nor_0.A
rlabel via1 1620 435 1620 435 1 L
rlabel via1 1640 -315 1640 -315 1 G
rlabel via1 1245 -315 1245 -315 1 E
<< end >>
