* Extracted by KLayout with GF180MCU LVS runset on : 03/10/2025 15:39

.SUBCKT gf180mcu_gp9t3v3__comp2_1 VSS A L E G VDD B
M$1 VDD B \$18 VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U PD=2.24U
M$2 G \$24 VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U PD=4.48U
M$3 VDD \$21 L VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U PD=2.24U
M$4 \$16 A VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U PD=4.48U
M$5 \$24 \$18 VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U
+ PD=2.24U
M$6 VDD A \$24 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U PD=4.48U
M$7 \$21 B VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U PD=2.24U
M$8 VDD \$16 \$21 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.459P PS=2.24U
+ PD=2.24U
M$9 \$36 \$16 VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.459P PS=2.24U
+ PD=2.24U
M$10 E A \$36 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U PD=4.48U
M$11 \$36 B VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.918P AD=0.459P PS=4.48U
+ PD=2.24U
M$12 E \$18 \$36 VDD pfet_03v3 L=0.3U W=1.7U AS=0.459P AD=0.918P PS=2.24U
+ PD=4.48U
M$13 VSS B \$18 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$14 G \$24 VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.2295P AD=0.459P PS=1.39U
+ PD=2.78U
M$15 \$32 \$18 \$24 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.102P PS=2.78U
+ PD=1.09U
M$16 VSS A \$32 VSS nfet_03v3 L=0.3U W=0.85U AS=0.102P AD=0.459P PS=1.09U
+ PD=2.78U
M$17 VSS \$21 L VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$18 \$16 A VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.2295P AD=0.459P PS=1.39U
+ PD=2.78U
M$19 E \$16 \$17 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$20 \$29 A E VSS nfet_03v3 L=0.3U W=0.85U AS=0.2295P AD=0.459P PS=1.39U
+ PD=2.78U
M$21 VSS B \$17 VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.2295P PS=2.78U
+ PD=1.39U
M$22 \$29 \$18 VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.2295P AD=0.459P PS=1.39U
+ PD=2.78U
M$23 \$31 B VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.459P AD=0.102P PS=2.78U
+ PD=1.09U
M$24 \$21 \$16 \$31 VSS nfet_03v3 L=0.3U W=0.85U AS=0.102P AD=0.459P PS=1.09U
+ PD=2.78U
.ENDS gf180mcu_gp9t3v3__comp2_1
