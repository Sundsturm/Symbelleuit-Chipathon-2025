magic
tech gf180mcuD
magscale 1 10
timestamp 1759424761
<< nwell >>
rect -13378 13441 -9260 14153
<< nmos >>
rect -12969 13139 -12909 13309
rect -12801 13139 -12741 13309
rect -12633 13139 -12573 13309
rect -12297 13139 -12237 13309
rect -12189 13139 -12129 13309
rect -11853 13139 -11793 13309
rect -11685 13139 -11625 13309
rect -11517 13139 -11457 13309
rect -11181 13139 -11121 13309
rect -11013 13139 -10953 13309
rect -10845 13139 -10785 13309
rect -10509 13139 -10449 13309
rect -10401 13139 -10341 13309
rect -10065 13139 -10005 13309
rect -9897 13139 -9837 13309
rect -9729 13139 -9669 13309
<< pmos >>
rect -12945 13531 -12885 13871
rect -12777 13531 -12717 13871
rect -12609 13531 -12549 13871
rect -12273 13531 -12213 13871
rect -12105 13531 -12045 13871
rect -11937 13531 -11877 13871
rect -11769 13531 -11709 13871
rect -11601 13531 -11541 13871
rect -11265 13531 -11205 13871
rect -11097 13531 -11037 13871
rect -10929 13531 -10869 13871
rect -10593 13531 -10533 13871
rect -10425 13531 -10365 13871
rect -10089 13531 -10029 13871
rect -9921 13531 -9861 13871
rect -9753 13531 -9693 13871
<< ndiff >>
rect -13077 13247 -12969 13309
rect -13077 13201 -13046 13247
rect -13000 13201 -12969 13247
rect -13077 13139 -12969 13201
rect -12909 13247 -12801 13309
rect -12909 13201 -12878 13247
rect -12832 13201 -12801 13247
rect -12909 13139 -12801 13201
rect -12741 13247 -12633 13309
rect -12741 13201 -12710 13247
rect -12664 13201 -12633 13247
rect -12741 13139 -12633 13201
rect -12573 13247 -12465 13309
rect -12573 13201 -12542 13247
rect -12496 13201 -12465 13247
rect -12573 13139 -12465 13201
rect -12405 13247 -12297 13309
rect -12405 13201 -12374 13247
rect -12328 13201 -12297 13247
rect -12405 13139 -12297 13201
rect -12237 13139 -12189 13309
rect -12129 13247 -12021 13309
rect -12129 13201 -12098 13247
rect -12052 13201 -12021 13247
rect -12129 13139 -12021 13201
rect -11961 13247 -11853 13309
rect -11961 13201 -11930 13247
rect -11884 13201 -11853 13247
rect -11961 13139 -11853 13201
rect -11793 13247 -11685 13309
rect -11793 13201 -11762 13247
rect -11716 13201 -11685 13247
rect -11793 13139 -11685 13201
rect -11625 13247 -11517 13309
rect -11625 13201 -11594 13247
rect -11548 13201 -11517 13247
rect -11625 13139 -11517 13201
rect -11457 13247 -11349 13309
rect -11457 13201 -11426 13247
rect -11380 13201 -11349 13247
rect -11457 13139 -11349 13201
rect -11289 13247 -11181 13309
rect -11289 13201 -11258 13247
rect -11212 13201 -11181 13247
rect -11289 13139 -11181 13201
rect -11121 13247 -11013 13309
rect -11121 13201 -11090 13247
rect -11044 13201 -11013 13247
rect -11121 13139 -11013 13201
rect -10953 13247 -10845 13309
rect -10953 13201 -10922 13247
rect -10876 13201 -10845 13247
rect -10953 13139 -10845 13201
rect -10785 13247 -10677 13309
rect -10785 13201 -10754 13247
rect -10708 13201 -10677 13247
rect -10785 13139 -10677 13201
rect -10617 13247 -10509 13309
rect -10617 13201 -10586 13247
rect -10540 13201 -10509 13247
rect -10617 13139 -10509 13201
rect -10449 13139 -10401 13309
rect -10341 13247 -10233 13309
rect -10341 13201 -10310 13247
rect -10264 13201 -10233 13247
rect -10341 13139 -10233 13201
rect -10173 13247 -10065 13309
rect -10173 13201 -10142 13247
rect -10096 13201 -10065 13247
rect -10173 13139 -10065 13201
rect -10005 13247 -9897 13309
rect -10005 13201 -9974 13247
rect -9928 13201 -9897 13247
rect -10005 13139 -9897 13201
rect -9837 13247 -9729 13309
rect -9837 13201 -9806 13247
rect -9760 13201 -9729 13247
rect -9837 13139 -9729 13201
rect -9669 13247 -9561 13309
rect -9669 13201 -9638 13247
rect -9592 13201 -9561 13247
rect -9669 13139 -9561 13201
<< pdiff >>
rect -13053 13818 -12945 13871
rect -13053 13584 -13022 13818
rect -12976 13584 -12945 13818
rect -13053 13531 -12945 13584
rect -12885 13818 -12777 13871
rect -12885 13584 -12854 13818
rect -12808 13584 -12777 13818
rect -12885 13531 -12777 13584
rect -12717 13818 -12609 13871
rect -12717 13584 -12686 13818
rect -12640 13584 -12609 13818
rect -12717 13531 -12609 13584
rect -12549 13818 -12441 13871
rect -12549 13584 -12518 13818
rect -12472 13584 -12441 13818
rect -12549 13531 -12441 13584
rect -12381 13818 -12273 13871
rect -12381 13584 -12350 13818
rect -12304 13584 -12273 13818
rect -12381 13531 -12273 13584
rect -12213 13818 -12105 13871
rect -12213 13584 -12182 13818
rect -12136 13584 -12105 13818
rect -12213 13531 -12105 13584
rect -12045 13818 -11937 13871
rect -12045 13584 -12014 13818
rect -11968 13584 -11937 13818
rect -12045 13531 -11937 13584
rect -11877 13818 -11769 13871
rect -11877 13584 -11846 13818
rect -11800 13584 -11769 13818
rect -11877 13531 -11769 13584
rect -11709 13818 -11601 13871
rect -11709 13584 -11678 13818
rect -11632 13584 -11601 13818
rect -11709 13531 -11601 13584
rect -11541 13818 -11433 13871
rect -11541 13584 -11510 13818
rect -11464 13584 -11433 13818
rect -11541 13531 -11433 13584
rect -11373 13818 -11265 13871
rect -11373 13584 -11342 13818
rect -11296 13584 -11265 13818
rect -11373 13531 -11265 13584
rect -11205 13818 -11097 13871
rect -11205 13584 -11174 13818
rect -11128 13584 -11097 13818
rect -11205 13531 -11097 13584
rect -11037 13818 -10929 13871
rect -11037 13584 -11006 13818
rect -10960 13584 -10929 13818
rect -11037 13531 -10929 13584
rect -10869 13818 -10761 13871
rect -10869 13584 -10838 13818
rect -10792 13584 -10761 13818
rect -10869 13531 -10761 13584
rect -10701 13818 -10593 13871
rect -10701 13584 -10670 13818
rect -10624 13584 -10593 13818
rect -10701 13531 -10593 13584
rect -10533 13818 -10425 13871
rect -10533 13584 -10502 13818
rect -10456 13584 -10425 13818
rect -10533 13531 -10425 13584
rect -10365 13818 -10257 13871
rect -10365 13584 -10334 13818
rect -10288 13584 -10257 13818
rect -10365 13531 -10257 13584
rect -10197 13818 -10089 13871
rect -10197 13584 -10166 13818
rect -10120 13584 -10089 13818
rect -10197 13531 -10089 13584
rect -10029 13818 -9921 13871
rect -10029 13584 -9998 13818
rect -9952 13584 -9921 13818
rect -10029 13531 -9921 13584
rect -9861 13818 -9753 13871
rect -9861 13584 -9830 13818
rect -9784 13584 -9753 13818
rect -9861 13531 -9753 13584
rect -9693 13818 -9585 13871
rect -9693 13584 -9662 13818
rect -9616 13584 -9585 13818
rect -9693 13531 -9585 13584
<< ndiffc >>
rect -13046 13201 -13000 13247
rect -12878 13201 -12832 13247
rect -12710 13201 -12664 13247
rect -12542 13201 -12496 13247
rect -12374 13201 -12328 13247
rect -12098 13201 -12052 13247
rect -11930 13201 -11884 13247
rect -11762 13201 -11716 13247
rect -11594 13201 -11548 13247
rect -11426 13201 -11380 13247
rect -11258 13201 -11212 13247
rect -11090 13201 -11044 13247
rect -10922 13201 -10876 13247
rect -10754 13201 -10708 13247
rect -10586 13201 -10540 13247
rect -10310 13201 -10264 13247
rect -10142 13201 -10096 13247
rect -9974 13201 -9928 13247
rect -9806 13201 -9760 13247
rect -9638 13201 -9592 13247
<< pdiffc >>
rect -13022 13584 -12976 13818
rect -12854 13584 -12808 13818
rect -12686 13584 -12640 13818
rect -12518 13584 -12472 13818
rect -12350 13584 -12304 13818
rect -12182 13584 -12136 13818
rect -12014 13584 -11968 13818
rect -11846 13584 -11800 13818
rect -11678 13584 -11632 13818
rect -11510 13584 -11464 13818
rect -11342 13584 -11296 13818
rect -11174 13584 -11128 13818
rect -11006 13584 -10960 13818
rect -10838 13584 -10792 13818
rect -10670 13584 -10624 13818
rect -10502 13584 -10456 13818
rect -10334 13584 -10288 13818
rect -10166 13584 -10120 13818
rect -9998 13584 -9952 13818
rect -9830 13584 -9784 13818
rect -9662 13584 -9616 13818
<< psubdiff >>
rect -13314 12955 -13164 12977
rect -13314 12909 -13262 12955
rect -13216 12909 -13164 12955
rect -13314 12887 -13164 12909
rect -13074 12955 -12924 12977
rect -13074 12909 -13022 12955
rect -12976 12909 -12924 12955
rect -13074 12887 -12924 12909
rect -12834 12955 -12684 12977
rect -12834 12909 -12782 12955
rect -12736 12909 -12684 12955
rect -12834 12887 -12684 12909
rect -12594 12955 -12444 12977
rect -12594 12909 -12542 12955
rect -12496 12909 -12444 12955
rect -12594 12887 -12444 12909
rect -12354 12955 -12204 12977
rect -12354 12909 -12302 12955
rect -12256 12909 -12204 12955
rect -12354 12887 -12204 12909
rect -12114 12955 -11964 12977
rect -12114 12909 -12062 12955
rect -12016 12909 -11964 12955
rect -12114 12887 -11964 12909
rect -11874 12955 -11724 12977
rect -11874 12909 -11822 12955
rect -11776 12909 -11724 12955
rect -11874 12887 -11724 12909
rect -11634 12955 -11484 12977
rect -11634 12909 -11582 12955
rect -11536 12909 -11484 12955
rect -11634 12887 -11484 12909
rect -11394 12955 -11244 12977
rect -11394 12909 -11342 12955
rect -11296 12909 -11244 12955
rect -11394 12887 -11244 12909
rect -11154 12955 -11004 12977
rect -11154 12909 -11102 12955
rect -11056 12909 -11004 12955
rect -11154 12887 -11004 12909
rect -10914 12955 -10764 12977
rect -10914 12909 -10862 12955
rect -10816 12909 -10764 12955
rect -10914 12887 -10764 12909
rect -10674 12955 -10524 12977
rect -10674 12909 -10622 12955
rect -10576 12909 -10524 12955
rect -10674 12887 -10524 12909
rect -10434 12955 -10284 12977
rect -10434 12909 -10382 12955
rect -10336 12909 -10284 12955
rect -10434 12887 -10284 12909
rect -10194 12955 -10044 12977
rect -10194 12909 -10142 12955
rect -10096 12909 -10044 12955
rect -10194 12887 -10044 12909
rect -9954 12955 -9804 12977
rect -9954 12909 -9902 12955
rect -9856 12909 -9804 12955
rect -9954 12887 -9804 12909
rect -9714 12955 -9564 12977
rect -9714 12909 -9662 12955
rect -9616 12909 -9564 12955
rect -9714 12887 -9564 12909
rect -9474 12955 -9324 12977
rect -9474 12909 -9422 12955
rect -9376 12909 -9324 12955
rect -9474 12887 -9324 12909
<< nsubdiff >>
rect -13314 14099 -13164 14121
rect -13314 14053 -13262 14099
rect -13216 14053 -13164 14099
rect -13314 14031 -13164 14053
rect -13074 14099 -12924 14121
rect -13074 14053 -13022 14099
rect -12976 14053 -12924 14099
rect -13074 14031 -12924 14053
rect -12834 14099 -12684 14121
rect -12834 14053 -12782 14099
rect -12736 14053 -12684 14099
rect -12834 14031 -12684 14053
rect -12594 14099 -12444 14121
rect -12594 14053 -12542 14099
rect -12496 14053 -12444 14099
rect -12594 14031 -12444 14053
rect -12354 14099 -12204 14121
rect -12354 14053 -12302 14099
rect -12256 14053 -12204 14099
rect -12354 14031 -12204 14053
rect -12114 14099 -11964 14121
rect -12114 14053 -12062 14099
rect -12016 14053 -11964 14099
rect -12114 14031 -11964 14053
rect -11874 14099 -11724 14121
rect -11874 14053 -11822 14099
rect -11776 14053 -11724 14099
rect -11874 14031 -11724 14053
rect -11634 14099 -11484 14121
rect -11634 14053 -11582 14099
rect -11536 14053 -11484 14099
rect -11634 14031 -11484 14053
rect -11394 14099 -11244 14121
rect -11394 14053 -11342 14099
rect -11296 14053 -11244 14099
rect -11394 14031 -11244 14053
rect -11154 14099 -11004 14121
rect -11154 14053 -11102 14099
rect -11056 14053 -11004 14099
rect -11154 14031 -11004 14053
rect -10914 14099 -10764 14121
rect -10914 14053 -10862 14099
rect -10816 14053 -10764 14099
rect -10914 14031 -10764 14053
rect -10674 14099 -10524 14121
rect -10674 14053 -10622 14099
rect -10576 14053 -10524 14099
rect -10674 14031 -10524 14053
rect -10434 14099 -10284 14121
rect -10434 14053 -10382 14099
rect -10336 14053 -10284 14099
rect -10434 14031 -10284 14053
rect -10194 14099 -10044 14121
rect -10194 14053 -10142 14099
rect -10096 14053 -10044 14099
rect -10194 14031 -10044 14053
rect -9954 14099 -9804 14121
rect -9954 14053 -9902 14099
rect -9856 14053 -9804 14099
rect -9954 14031 -9804 14053
rect -9714 14099 -9564 14121
rect -9714 14053 -9662 14099
rect -9616 14053 -9564 14099
rect -9714 14031 -9564 14053
rect -9474 14099 -9324 14121
rect -9474 14053 -9422 14099
rect -9376 14053 -9324 14099
rect -9474 14031 -9324 14053
<< psubdiffcont >>
rect -13262 12909 -13216 12955
rect -13022 12909 -12976 12955
rect -12782 12909 -12736 12955
rect -12542 12909 -12496 12955
rect -12302 12909 -12256 12955
rect -12062 12909 -12016 12955
rect -11822 12909 -11776 12955
rect -11582 12909 -11536 12955
rect -11342 12909 -11296 12955
rect -11102 12909 -11056 12955
rect -10862 12909 -10816 12955
rect -10622 12909 -10576 12955
rect -10382 12909 -10336 12955
rect -10142 12909 -10096 12955
rect -9902 12909 -9856 12955
rect -9662 12909 -9616 12955
rect -9422 12909 -9376 12955
<< nsubdiffcont >>
rect -13262 14053 -13216 14099
rect -13022 14053 -12976 14099
rect -12782 14053 -12736 14099
rect -12542 14053 -12496 14099
rect -12302 14053 -12256 14099
rect -12062 14053 -12016 14099
rect -11822 14053 -11776 14099
rect -11582 14053 -11536 14099
rect -11342 14053 -11296 14099
rect -11102 14053 -11056 14099
rect -10862 14053 -10816 14099
rect -10622 14053 -10576 14099
rect -10382 14053 -10336 14099
rect -10142 14053 -10096 14099
rect -9902 14053 -9856 14099
rect -9662 14053 -9616 14099
rect -9422 14053 -9376 14099
<< polysilicon >>
rect -12273 13969 -10029 14009
rect -12945 13871 -12885 13921
rect -12777 13871 -12717 13921
rect -12609 13871 -12549 13921
rect -12273 13871 -12213 13969
rect -12105 13871 -12045 13921
rect -11937 13871 -11877 13921
rect -11769 13871 -11709 13921
rect -11601 13871 -11541 13921
rect -11265 13871 -11205 13969
rect -11097 13871 -11037 13921
rect -10929 13871 -10869 13921
rect -10593 13871 -10533 13921
rect -10425 13871 -10365 13921
rect -10089 13871 -10029 13969
rect -9921 13871 -9861 13921
rect -9753 13871 -9693 13921
rect -12945 13511 -12885 13531
rect -12777 13511 -12717 13531
rect -12945 13471 -12717 13511
rect -12801 13455 -12717 13471
rect -12801 13409 -12782 13455
rect -12736 13409 -12717 13455
rect -12801 13369 -12717 13409
rect -12609 13369 -12549 13531
rect -12273 13511 -12213 13531
rect -12297 13471 -12213 13511
rect -12337 13447 -12237 13471
rect -12337 13401 -12311 13447
rect -12265 13401 -12237 13447
rect -12337 13371 -12237 13401
rect -12105 13462 -12045 13531
rect -11937 13462 -11877 13531
rect -11769 13511 -11709 13531
rect -11601 13511 -11541 13531
rect -11265 13511 -11205 13531
rect -11097 13511 -11037 13531
rect -11769 13471 -11457 13511
rect -12105 13443 -11877 13462
rect -12105 13397 -12014 13443
rect -11968 13397 -11877 13443
rect -12105 13377 -11877 13397
rect -12969 13329 -12741 13369
rect -12969 13309 -12909 13329
rect -12801 13309 -12741 13329
rect -12633 13329 -12549 13369
rect -12633 13309 -12573 13329
rect -12297 13309 -12237 13371
rect -12189 13337 -11793 13377
rect -11517 13369 -11457 13471
rect -12189 13309 -12129 13337
rect -11853 13309 -11793 13337
rect -11685 13329 -11457 13369
rect -11265 13471 -11037 13511
rect -10929 13511 -10869 13531
rect -10593 13511 -10533 13531
rect -10929 13471 -10533 13511
rect -10425 13511 -10365 13531
rect -10425 13471 -10341 13511
rect -11265 13369 -11205 13471
rect -10654 13441 -10554 13471
rect -10654 13395 -10627 13441
rect -10581 13395 -10554 13441
rect -10654 13369 -10554 13395
rect -10401 13447 -10241 13471
rect -10401 13401 -10315 13447
rect -10269 13401 -10241 13447
rect -10401 13371 -10241 13401
rect -10089 13377 -10029 13531
rect -9921 13511 -9861 13531
rect -9753 13511 -9693 13531
rect -9921 13471 -9693 13511
rect -9921 13455 -9837 13471
rect -9921 13409 -9902 13455
rect -9856 13409 -9837 13455
rect -11265 13329 -11121 13369
rect -11685 13309 -11625 13329
rect -11517 13309 -11457 13329
rect -11181 13309 -11121 13329
rect -11013 13329 -10449 13369
rect -11013 13309 -10953 13329
rect -10845 13309 -10785 13329
rect -10509 13309 -10449 13329
rect -10401 13309 -10341 13371
rect -10089 13337 -10005 13377
rect -9921 13369 -9837 13409
rect -10065 13309 -10005 13337
rect -9897 13329 -9669 13369
rect -9897 13309 -9837 13329
rect -9729 13309 -9669 13329
rect -12969 13089 -12909 13139
rect -12801 13089 -12741 13139
rect -12633 13041 -12573 13139
rect -12297 13089 -12237 13139
rect -12189 13089 -12129 13139
rect -11853 13089 -11793 13139
rect -11685 13089 -11625 13139
rect -11517 13041 -11457 13139
rect -11181 13089 -11121 13139
rect -11013 13089 -10953 13139
rect -10845 13089 -10785 13139
rect -10509 13089 -10449 13139
rect -10401 13041 -10341 13139
rect -10065 13089 -10005 13139
rect -9897 13089 -9837 13139
rect -9729 13089 -9669 13139
rect -12633 13001 -10341 13041
<< polycontact >>
rect -12782 13409 -12736 13455
rect -12311 13401 -12265 13447
rect -12014 13397 -11968 13443
rect -10627 13395 -10581 13441
rect -10315 13401 -10269 13447
rect -9902 13409 -9856 13455
<< metal1 >>
rect -13378 14099 -9260 14153
rect -13378 14053 -13262 14099
rect -13216 14053 -13022 14099
rect -12976 14053 -12782 14099
rect -12736 14053 -12542 14099
rect -12496 14053 -12302 14099
rect -12256 14053 -12062 14099
rect -12016 14053 -11822 14099
rect -11776 14053 -11582 14099
rect -11536 14053 -11342 14099
rect -11296 14053 -11102 14099
rect -11056 14053 -10862 14099
rect -10816 14053 -10622 14099
rect -10576 14053 -10382 14099
rect -10336 14053 -10142 14099
rect -10096 14053 -9902 14099
rect -9856 14053 -9662 14099
rect -9616 14053 -9422 14099
rect -9376 14053 -9260 14099
rect -13378 14013 -9260 14053
rect -13025 13818 -12973 14013
rect -13025 13584 -13022 13818
rect -12976 13584 -12973 13818
rect -13025 13531 -12973 13584
rect -12858 13818 -12806 13871
rect -12858 13584 -12854 13818
rect -12808 13584 -12806 13818
rect -12858 13583 -12806 13584
rect -12911 13531 -12806 13583
rect -12689 13818 -12637 14013
rect -12689 13584 -12686 13818
rect -12640 13584 -12637 13818
rect -12689 13531 -12637 13584
rect -12522 13818 -12470 13874
rect -12522 13584 -12518 13818
rect -12472 13584 -12470 13818
rect -12911 13475 -12859 13531
rect -12522 13513 -12470 13584
rect -12353 13818 -12301 14013
rect -12353 13584 -12350 13818
rect -12304 13584 -12301 13818
rect -12353 13559 -12301 13584
rect -12185 13818 -12133 13871
rect -12185 13584 -12182 13818
rect -12136 13584 -12133 13818
rect -12960 13458 -12859 13475
rect -12960 13406 -12936 13458
rect -12884 13406 -12859 13458
rect -12960 13379 -12859 13406
rect -12801 13458 -12717 13475
rect -12801 13406 -12785 13458
rect -12733 13406 -12717 13458
rect -12801 13379 -12717 13406
rect -12546 13471 -12470 13513
rect -12546 13419 -12535 13471
rect -12483 13419 -12470 13471
rect -12909 13309 -12859 13379
rect -12546 13337 -12470 13419
rect -12337 13485 -12237 13511
rect -12337 13433 -12321 13485
rect -12269 13447 -12237 13485
rect -12337 13401 -12311 13433
rect -12265 13401 -12237 13447
rect -12337 13371 -12237 13401
rect -13049 13247 -12997 13309
rect -12909 13257 -12829 13309
rect -13049 13201 -13046 13247
rect -13000 13201 -12997 13247
rect -13049 13023 -12997 13201
rect -12881 13247 -12829 13257
rect -12881 13201 -12878 13247
rect -12832 13201 -12829 13247
rect -12881 13134 -12829 13201
rect -12713 13247 -12661 13309
rect -12713 13201 -12710 13247
rect -12664 13201 -12661 13247
rect -12713 13023 -12661 13201
rect -12546 13247 -12494 13337
rect -12185 13309 -12133 13584
rect -12017 13818 -11965 14013
rect -12017 13584 -12014 13818
rect -11968 13584 -11965 13818
rect -12017 13531 -11965 13584
rect -11849 13818 -11797 13878
rect -11849 13584 -11846 13818
rect -11800 13584 -11797 13818
rect -11849 13512 -11797 13584
rect -11709 13818 -11601 13871
rect -11709 13779 -11678 13818
rect -11632 13779 -11601 13818
rect -11709 13623 -11681 13779
rect -11629 13623 -11601 13779
rect -11709 13584 -11678 13623
rect -11632 13584 -11601 13623
rect -11709 13560 -11601 13584
rect -11513 13818 -11461 13871
rect -11513 13584 -11510 13818
rect -11464 13584 -11461 13818
rect -11513 13512 -11461 13584
rect -11345 13818 -11293 13871
rect -11345 13584 -11342 13818
rect -11296 13584 -11293 13818
rect -11345 13512 -11293 13584
rect -11177 13818 -11125 14013
rect -11177 13584 -11174 13818
rect -11128 13584 -11125 13818
rect -11177 13560 -11125 13584
rect -11009 13818 -10957 13871
rect -11009 13584 -11006 13818
rect -10960 13584 -10957 13818
rect -11009 13512 -10957 13584
rect -10869 13818 -10761 13871
rect -10869 13779 -10838 13818
rect -10792 13779 -10761 13818
rect -10869 13623 -10841 13779
rect -10789 13623 -10761 13779
rect -10869 13584 -10838 13623
rect -10792 13584 -10761 13623
rect -10869 13560 -10761 13584
rect -10673 13818 -10621 14013
rect -10673 13584 -10670 13818
rect -10624 13584 -10621 13818
rect -10673 13531 -10621 13584
rect -10505 13818 -10453 13871
rect -10505 13584 -10502 13818
rect -10456 13584 -10453 13818
rect -12045 13446 -11937 13462
rect -11849 13460 -10957 13512
rect -12045 13394 -12017 13446
rect -11965 13394 -11937 13446
rect -10654 13444 -10554 13463
rect -12045 13377 -11937 13394
rect -11597 13357 -10873 13409
rect -10654 13392 -10630 13444
rect -10578 13392 -10554 13444
rect -10654 13377 -10554 13392
rect -12546 13201 -12542 13247
rect -12496 13201 -12494 13247
rect -12546 13139 -12494 13201
rect -12377 13247 -12325 13309
rect -12377 13201 -12374 13247
rect -12328 13201 -12325 13247
rect -12377 13023 -12325 13201
rect -12189 13247 -12021 13309
rect -12189 13214 -12098 13247
rect -12052 13214 -12021 13247
rect -12189 13162 -12101 13214
rect -12049 13162 -12021 13214
rect -12189 13139 -12021 13162
rect -11933 13247 -11881 13309
rect -11933 13201 -11930 13247
rect -11884 13201 -11881 13247
rect -11933 13123 -11881 13201
rect -11793 13249 -11685 13278
rect -11793 13197 -11765 13249
rect -11713 13197 -11685 13249
rect -11793 13170 -11685 13197
rect -11597 13247 -11545 13357
rect -11597 13201 -11594 13247
rect -11548 13201 -11545 13247
rect -11597 13171 -11545 13201
rect -11457 13249 -11349 13278
rect -11457 13197 -11429 13249
rect -11377 13197 -11349 13249
rect -11457 13170 -11349 13197
rect -11261 13247 -11209 13309
rect -11261 13201 -11258 13247
rect -11212 13201 -11209 13247
rect -11261 13123 -11209 13201
rect -11934 13071 -11209 13123
rect -11093 13247 -11041 13309
rect -11093 13201 -11090 13247
rect -11044 13201 -11041 13247
rect -11093 13023 -11041 13201
rect -10925 13247 -10873 13357
rect -10505 13309 -10453 13584
rect -10337 13818 -10285 14013
rect -10337 13584 -10334 13818
rect -10288 13584 -10285 13818
rect -10337 13559 -10285 13584
rect -10169 13818 -10117 13874
rect -10169 13584 -10166 13818
rect -10120 13584 -10117 13818
rect -10169 13513 -10117 13584
rect -10001 13818 -9949 14013
rect -10001 13584 -9998 13818
rect -9952 13584 -9949 13818
rect -10001 13531 -9949 13584
rect -9833 13818 -9781 13871
rect -9833 13584 -9830 13818
rect -9784 13584 -9781 13818
rect -9833 13583 -9781 13584
rect -9665 13818 -9613 14013
rect -9665 13584 -9662 13818
rect -9616 13584 -9613 13818
rect -9833 13531 -9729 13583
rect -9665 13531 -9613 13584
rect -10341 13485 -10241 13511
rect -10341 13433 -10325 13485
rect -10273 13447 -10241 13485
rect -10341 13401 -10315 13433
rect -10269 13401 -10241 13447
rect -10341 13371 -10241 13401
rect -10169 13471 -10093 13513
rect -9781 13480 -9729 13531
rect -10169 13419 -10156 13471
rect -10104 13419 -10093 13471
rect -10169 13377 -10093 13419
rect -9921 13458 -9837 13480
rect -9921 13406 -9905 13458
rect -9853 13406 -9837 13458
rect -9921 13379 -9837 13406
rect -9781 13458 -9678 13480
rect -9781 13406 -9753 13458
rect -9701 13406 -9678 13458
rect -9781 13379 -9678 13406
rect -10925 13201 -10922 13247
rect -10876 13201 -10873 13247
rect -10925 13139 -10873 13201
rect -10757 13247 -10705 13309
rect -10757 13201 -10754 13247
rect -10708 13201 -10705 13247
rect -10757 13023 -10705 13201
rect -10617 13247 -10449 13309
rect -10617 13218 -10586 13247
rect -10540 13218 -10449 13247
rect -10617 13166 -10589 13218
rect -10537 13166 -10449 13218
rect -10617 13139 -10449 13166
rect -10313 13247 -10261 13309
rect -10313 13201 -10310 13247
rect -10264 13201 -10261 13247
rect -10313 13023 -10261 13201
rect -10145 13247 -10093 13377
rect -9781 13309 -9729 13379
rect -10145 13201 -10142 13247
rect -10096 13201 -10093 13247
rect -10145 13139 -10093 13201
rect -9977 13247 -9925 13309
rect -9977 13201 -9974 13247
rect -9928 13201 -9925 13247
rect -9977 13023 -9925 13201
rect -9809 13257 -9729 13309
rect -9809 13247 -9757 13257
rect -9809 13201 -9806 13247
rect -9760 13201 -9757 13247
rect -9809 13140 -9757 13201
rect -9641 13247 -9589 13309
rect -9641 13201 -9638 13247
rect -9592 13201 -9589 13247
rect -9641 13023 -9589 13201
rect -13378 12955 -9260 13023
rect -13378 12909 -13262 12955
rect -13216 12909 -13022 12955
rect -12976 12909 -12782 12955
rect -12736 12909 -12542 12955
rect -12496 12909 -12302 12955
rect -12256 12909 -12062 12955
rect -12016 12909 -11822 12955
rect -11776 12909 -11582 12955
rect -11536 12909 -11342 12955
rect -11296 12909 -11102 12955
rect -11056 12909 -10862 12955
rect -10816 12909 -10622 12955
rect -10576 12909 -10382 12955
rect -10336 12909 -10142 12955
rect -10096 12909 -9902 12955
rect -9856 12909 -9662 12955
rect -9616 12909 -9422 12955
rect -9376 12909 -9260 12955
rect -13378 12883 -9260 12909
<< via1 >>
rect -12936 13406 -12884 13458
rect -12785 13455 -12733 13458
rect -12785 13409 -12782 13455
rect -12782 13409 -12736 13455
rect -12736 13409 -12733 13455
rect -12785 13406 -12733 13409
rect -12535 13419 -12483 13471
rect -12321 13447 -12269 13485
rect -12321 13433 -12311 13447
rect -12311 13433 -12269 13447
rect -11681 13623 -11678 13779
rect -11678 13623 -11632 13779
rect -11632 13623 -11629 13779
rect -10841 13623 -10838 13779
rect -10838 13623 -10792 13779
rect -10792 13623 -10789 13779
rect -12017 13443 -11965 13446
rect -12017 13397 -12014 13443
rect -12014 13397 -11968 13443
rect -11968 13397 -11965 13443
rect -12017 13394 -11965 13397
rect -10630 13441 -10578 13444
rect -10630 13395 -10627 13441
rect -10627 13395 -10581 13441
rect -10581 13395 -10578 13441
rect -10630 13392 -10578 13395
rect -12101 13201 -12098 13214
rect -12098 13201 -12052 13214
rect -12052 13201 -12049 13214
rect -12101 13162 -12049 13201
rect -11765 13247 -11713 13249
rect -11765 13201 -11762 13247
rect -11762 13201 -11716 13247
rect -11716 13201 -11713 13247
rect -11765 13197 -11713 13201
rect -11429 13247 -11377 13249
rect -11429 13201 -11426 13247
rect -11426 13201 -11380 13247
rect -11380 13201 -11377 13247
rect -11429 13197 -11377 13201
rect -10325 13447 -10273 13485
rect -10325 13433 -10315 13447
rect -10315 13433 -10273 13447
rect -10156 13419 -10104 13471
rect -9905 13455 -9853 13458
rect -9905 13409 -9902 13455
rect -9902 13409 -9856 13455
rect -9856 13409 -9853 13455
rect -9905 13406 -9853 13409
rect -9753 13406 -9701 13458
rect -10589 13201 -10586 13218
rect -10586 13201 -10540 13218
rect -10540 13201 -10537 13218
rect -10589 13166 -10537 13201
<< metal2 >>
rect -11709 13779 -11601 13871
rect -11709 13623 -11681 13779
rect -11629 13730 -11601 13779
rect -10869 13779 -10761 13871
rect -10869 13730 -10841 13779
rect -11629 13670 -10841 13730
rect -11629 13623 -11601 13670
rect -12960 13458 -12859 13475
rect -12960 13406 -12936 13458
rect -12884 13406 -12859 13458
rect -12960 13379 -12859 13406
rect -12801 13458 -12717 13503
rect -12801 13406 -12785 13458
rect -12733 13406 -12717 13458
rect -12546 13471 -12470 13513
rect -12546 13429 -12535 13471
rect -12801 13379 -12717 13406
rect -12537 13419 -12535 13429
rect -12483 13429 -12470 13471
rect -12337 13485 -12253 13511
rect -12337 13433 -12321 13485
rect -12269 13433 -12253 13485
rect -12483 13419 -12477 13429
rect -12801 13153 -12741 13379
rect -12537 13357 -12477 13419
rect -12337 13417 -12253 13433
rect -12045 13446 -11937 13462
rect -12045 13394 -12017 13446
rect -11965 13394 -11937 13446
rect -12045 13377 -11937 13394
rect -12045 13357 -11985 13377
rect -12537 13297 -11985 13357
rect -11709 13278 -11601 13623
rect -10869 13623 -10841 13670
rect -10789 13623 -10761 13779
rect -10869 13560 -10761 13623
rect -10341 13485 -10257 13511
rect -10654 13444 -10554 13471
rect -10654 13392 -10630 13444
rect -10578 13392 -10554 13444
rect -10341 13433 -10325 13485
rect -10273 13433 -10257 13485
rect -10341 13417 -10257 13433
rect -10169 13471 -10093 13513
rect -9897 13480 -9837 13503
rect -10169 13419 -10156 13471
rect -10104 13419 -10093 13471
rect -10654 13377 -10554 13392
rect -10614 13357 -10554 13377
rect -10169 13377 -10093 13419
rect -9921 13458 -9837 13480
rect -9921 13406 -9905 13458
rect -9853 13406 -9837 13458
rect -9921 13379 -9837 13406
rect -9781 13458 -9678 13480
rect -9781 13406 -9753 13458
rect -9701 13406 -9678 13458
rect -9781 13379 -9678 13406
rect -10169 13357 -10109 13377
rect -10614 13297 -10109 13357
rect -11793 13249 -11349 13278
rect -12129 13214 -12021 13236
rect -12129 13162 -12101 13214
rect -12049 13162 -12021 13214
rect -11793 13197 -11765 13249
rect -11713 13197 -11429 13249
rect -11377 13197 -11349 13249
rect -11793 13170 -11349 13197
rect -10617 13218 -10449 13237
rect -12129 13153 -12021 13162
rect -12801 13093 -12021 13153
rect -10617 13166 -10589 13218
rect -10537 13199 -10449 13218
rect -9897 13199 -9837 13379
rect -10537 13166 -9837 13199
rect -10617 13139 -9837 13166
<< labels >>
flabel metal2 s -12288 13495 -12288 13495 2 FreeSans 448 0 0 0 B
port 1 nsew
flabel metal2 s -10296 13477 -10296 13477 2 FreeSans 448 0 0 0 A
port 2 nsew
flabel metal2 s -9764 13388 -9764 13388 2 FreeSans 700 0 0 0 G
port 3 nsew
flabel metal2 s -12918 13426 -12918 13426 2 FreeSans 700 0 0 0 L
port 4 nsew
flabel metal2 s -11643 13378 -11643 13378 2 FreeSans 700 0 0 0 E
port 5 nsew
flabel metal1 s -10244 14085 -10244 14085 2 FreeSans 576 0 0 0 VDD
port 6 nsew
flabel metal1 s -10244 12936 -10244 12936 2 FreeSans 576 0 0 0 VSS
port 7 nsew
<< properties >>
string path -62.535 67.145 -62.535 66.635 -60.075 66.635 -60.075 67.160 
<< end >>
